//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9.03 Education (64-bit)
//Part Number: GW1NR-LV9QN88PC6/I5
//Device: GW1NR-9
//Device Version: C
//Created Time: Sun Oct 13 20:10:48 2024

module Gowin_pROM (dout, clk, oce, ce, reset, ad);

output [1:0] dout;
input clk;
input oce;
input ce;
input reset;
input [17:0] ad;

wire lut_f_0;
wire lut_f_1;
wire lut_f_2;
wire lut_f_3;
wire lut_f_4;
wire lut_f_5;
wire lut_f_6;
wire lut_f_7;
wire lut_f_8;
wire lut_f_9;
wire lut_f_10;
wire lut_f_11;
wire lut_f_12;
wire lut_f_13;
wire lut_f_14;
wire lut_f_15;
wire lut_f_16;
wire lut_f_17;
wire lut_f_18;
wire lut_f_19;
wire [30:0] prom_inst_0_dout_w;
wire [0:0] prom_inst_0_dout;
wire [30:0] prom_inst_1_dout_w;
wire [0:0] prom_inst_1_dout;
wire [30:0] prom_inst_2_dout_w;
wire [0:0] prom_inst_2_dout;
wire [30:0] prom_inst_3_dout_w;
wire [0:0] prom_inst_3_dout;
wire [30:0] prom_inst_4_dout_w;
wire [0:0] prom_inst_4_dout;
wire [30:0] prom_inst_5_dout_w;
wire [0:0] prom_inst_5_dout;
wire [30:0] prom_inst_6_dout_w;
wire [0:0] prom_inst_6_dout;
wire [30:0] prom_inst_7_dout_w;
wire [0:0] prom_inst_7_dout;
wire [30:0] prom_inst_8_dout_w;
wire [1:1] prom_inst_8_dout;
wire [30:0] prom_inst_9_dout_w;
wire [1:1] prom_inst_9_dout;
wire [30:0] prom_inst_10_dout_w;
wire [1:1] prom_inst_10_dout;
wire [30:0] prom_inst_11_dout_w;
wire [1:1] prom_inst_11_dout;
wire [30:0] prom_inst_12_dout_w;
wire [1:1] prom_inst_12_dout;
wire [30:0] prom_inst_13_dout_w;
wire [1:1] prom_inst_13_dout;
wire [30:0] prom_inst_14_dout_w;
wire [1:1] prom_inst_14_dout;
wire [30:0] prom_inst_15_dout_w;
wire [1:1] prom_inst_15_dout;
wire [30:0] prom_inst_16_dout_w;
wire [0:0] prom_inst_16_dout;
wire [30:0] prom_inst_17_dout_w;
wire [1:1] prom_inst_17_dout;
wire [29:0] prom_inst_18_dout_w;
wire [1:0] prom_inst_18_dout;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire dff_q_3;
wire mux_o_10;
wire mux_o_11;
wire mux_o_12;
wire mux_o_13;
wire mux_o_14;
wire mux_o_15;
wire mux_o_16;
wire mux_o_18;
wire mux_o_31;
wire mux_o_32;
wire mux_o_33;
wire mux_o_34;
wire mux_o_35;
wire mux_o_36;
wire mux_o_37;
wire mux_o_39;
wire gw_gnd;

assign gw_gnd = 1'b0;

LUT4 lut_inst_0 (
  .F(lut_f_0),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17])
);
defparam lut_inst_0.INIT = 16'h0001;
LUT2 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(lut_f_0)
);
defparam lut_inst_1.INIT = 4'h8;
LUT4 lut_inst_2 (
  .F(lut_f_2),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17])
);
defparam lut_inst_2.INIT = 16'h0002;
LUT2 lut_inst_3 (
  .F(lut_f_3),
  .I0(ce),
  .I1(lut_f_2)
);
defparam lut_inst_3.INIT = 4'h8;
LUT4 lut_inst_4 (
  .F(lut_f_4),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17])
);
defparam lut_inst_4.INIT = 16'h0004;
LUT2 lut_inst_5 (
  .F(lut_f_5),
  .I0(ce),
  .I1(lut_f_4)
);
defparam lut_inst_5.INIT = 4'h8;
LUT4 lut_inst_6 (
  .F(lut_f_6),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17])
);
defparam lut_inst_6.INIT = 16'h0008;
LUT2 lut_inst_7 (
  .F(lut_f_7),
  .I0(ce),
  .I1(lut_f_6)
);
defparam lut_inst_7.INIT = 4'h8;
LUT4 lut_inst_8 (
  .F(lut_f_8),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17])
);
defparam lut_inst_8.INIT = 16'h0010;
LUT2 lut_inst_9 (
  .F(lut_f_9),
  .I0(ce),
  .I1(lut_f_8)
);
defparam lut_inst_9.INIT = 4'h8;
LUT4 lut_inst_10 (
  .F(lut_f_10),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17])
);
defparam lut_inst_10.INIT = 16'h0020;
LUT2 lut_inst_11 (
  .F(lut_f_11),
  .I0(ce),
  .I1(lut_f_10)
);
defparam lut_inst_11.INIT = 4'h8;
LUT4 lut_inst_12 (
  .F(lut_f_12),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17])
);
defparam lut_inst_12.INIT = 16'h0040;
LUT2 lut_inst_13 (
  .F(lut_f_13),
  .I0(ce),
  .I1(lut_f_12)
);
defparam lut_inst_13.INIT = 4'h8;
LUT4 lut_inst_14 (
  .F(lut_f_14),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17])
);
defparam lut_inst_14.INIT = 16'h0080;
LUT2 lut_inst_15 (
  .F(lut_f_15),
  .I0(ce),
  .I1(lut_f_14)
);
defparam lut_inst_15.INIT = 4'h8;
LUT4 lut_inst_16 (
  .F(lut_f_16),
  .I0(ad[14]),
  .I1(ad[15]),
  .I2(ad[16]),
  .I3(ad[17])
);
defparam lut_inst_16.INIT = 16'h0100;
LUT2 lut_inst_17 (
  .F(lut_f_17),
  .I0(ce),
  .I1(lut_f_16)
);
defparam lut_inst_17.INIT = 4'h8;
LUT5 lut_inst_18 (
  .F(lut_f_18),
  .I0(ad[13]),
  .I1(ad[14]),
  .I2(ad[15]),
  .I3(ad[16]),
  .I4(ad[17])
);
defparam lut_inst_18.INIT = 32'h00040000;
LUT2 lut_inst_19 (
  .F(lut_f_19),
  .I0(ce),
  .I1(lut_f_18)
);
defparam lut_inst_19.INIT = 4'h8;
pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],prom_inst_0_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[30:0],prom_inst_1_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 1;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_39 = 256'h0000000000000000000000002000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3F = 256'h0000000004000000000000000000000000000000000000000000000000000000;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[30:0],prom_inst_2_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_5),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 1;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000800000;
defparam prom_inst_2.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_09 = 256'h0000010000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000001000000000000000000000;
defparam prom_inst_2.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_12 = 256'h0000000000000000000000000002000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_13 = 256'h0000200000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_1A = 256'h0000000000000000000000000000400000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000020000000000000000000;
defparam prom_inst_2.INIT_RAM_1C = 256'h0000000000000000000200000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_20 = 256'h0000000000000800000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_21 = 256'h0000000000000000000000000000040000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_22 = 256'h0010000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_27 = 256'h0000000000000080000000000000000000000000000000000000000000000100;
defparam prom_inst_2.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000080000000000000;
defparam prom_inst_2.INIT_RAM_2A = 256'h0080000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000100;
defparam prom_inst_2.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000010000000000000;
defparam prom_inst_2.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000008000000000000000000;
defparam prom_inst_2.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_37 = 256'h0000000000000000000000000000000000020000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_38 = 256'h0000000000000000000000000000400000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_39 = 256'h000000000000000000000000000000000000000000000000C000000000000000;
defparam prom_inst_2.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3B = 256'h0000000000000000200000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000001;
defparam prom_inst_2.INIT_RAM_3D = 256'h0000000000000000200000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3E = 256'h0000000000000004000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[30:0],prom_inst_3_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_7),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 1;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000200000000000;
defparam prom_inst_3.INIT_RAM_01 = 256'h0400000000000000000000000000000000000000000400000000000000000000;
defparam prom_inst_3.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000080000000000000000;
defparam prom_inst_3.INIT_RAM_03 = 256'h0400000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000020;
defparam prom_inst_3.INIT_RAM_06 = 256'h0000000000000000000000000000000000000400000000000000000000000000;
defparam prom_inst_3.INIT_RAM_07 = 256'h0000000000000000010000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_08 = 256'h0000000000000000000000000000004000000100000000000080000000000000;
defparam prom_inst_3.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000001000000000000000000;
defparam prom_inst_3.INIT_RAM_0C = 256'h0000000000000000000000800000000000000000000000000000000000800000;
defparam prom_inst_3.INIT_RAM_0D = 256'h0020000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0E = 256'h0000000000000200000000200000000000100000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_11 = 256'h0000000000000000000000000000080000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_12 = 256'h0000001000000000000000000000000000000000040000000000000000000000;
defparam prom_inst_3.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_14 = 256'h0000000400000000000200000000000000000000000000000004000000000000;
defparam prom_inst_3.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000001000;
defparam prom_inst_3.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_17 = 256'h0000000000004000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_18 = 256'h0000000000004000000000002000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000200000000;
defparam prom_inst_3.INIT_RAM_1A = 256'h0000400000000000000000000000000000008000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000080000000;
defparam prom_inst_3.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000020000;
defparam prom_inst_3.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000020000;
defparam prom_inst_3.INIT_RAM_20 = 256'h0000000000000000000010000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_21 = 256'h0000000000000000000000000000000000000800000000000000000000000000;
defparam prom_inst_3.INIT_RAM_22 = 256'h0000080000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000020000100000;
defparam prom_inst_3.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000200000;
defparam prom_inst_3.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000010000000000;
defparam prom_inst_3.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_2B = 256'h0000000000000000000000000000000000000040008000000000000000000000;
defparam prom_inst_3.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_2D = 256'h0000008000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_2E = 256'h0000010000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_2F = 256'h0000000000000000000000000040000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_30 = 256'h0000020000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_31 = 256'h0000000000100000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000001000000000000000000000;
defparam prom_inst_3.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000040000000000;
defparam prom_inst_3.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000080000000000;
defparam prom_inst_3.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000100000000000;
defparam prom_inst_3.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000020000;
defparam prom_inst_3.INIT_RAM_39 = 256'h0000000000000000000000000002000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3B = 256'h0000000000000000000000000000000000004000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3C = 256'h0000000040000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3D = 256'h0000000040000000000000000000000000008000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3E = 256'h0000000180000000000000000000000000000000C00040000000000000000000;
defparam prom_inst_3.INIT_RAM_3F = 256'h000000020000400000000000C0000000000000000000000000000000E0000000;

pROM prom_inst_4 (
    .DO({prom_inst_4_dout_w[30:0],prom_inst_4_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_9),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_4.READ_MODE = 1'b0;
defparam prom_inst_4.BIT_WIDTH = 1;
defparam prom_inst_4.RESET_MODE = "SYNC";
defparam prom_inst_4.INIT_RAM_00 = 256'h00000001E0000000000000000000000000000000E00000000000000380000000;
defparam prom_inst_4.INIT_RAM_01 = 256'h000000000000000000020001F000000000000003C00000000000000020000000;
defparam prom_inst_4.INIT_RAM_02 = 256'h00000003F800000000000007C0000000000000000000000000000003F0001000;
defparam prom_inst_4.INIT_RAM_03 = 256'h00000007E0000000000400000000000000000003F00000000000000008000000;
defparam prom_inst_4.INIT_RAM_04 = 256'h000000000000000000080007F8000000000000000000000000000003F8000000;
defparam prom_inst_4.INIT_RAM_05 = 256'h0000000FF8000000000000000000000000000007FC0000000000000FF0000000;
defparam prom_inst_4.INIT_RAM_06 = 256'h000000000000000000000007FC0000000000001FF80000000000001000000800;
defparam prom_inst_4.INIT_RAM_07 = 256'h0000000FFE0000000000001FF800000000000000000000000010000FFC000000;
defparam prom_inst_4.INIT_RAM_08 = 256'h0000003FFC00000000000000000004000000001FFC0000000000000000000000;
defparam prom_inst_4.INIT_RAM_09 = 256'h00000000000000000000001FFE00000000000000000000000000001FFE000000;
defparam prom_inst_4.INIT_RAM_0A = 256'h0000003FFF00000000200000000000000000001FFF0000000000003FFC000000;
defparam prom_inst_4.INIT_RAM_0B = 256'h00000000008000000000003FFF8000000000007FFE0000000000000000000000;
defparam prom_inst_4.INIT_RAM_0C = 256'h0000003FFF800000000000FFFE00000000400000000000000000003FFF000000;
defparam prom_inst_4.INIT_RAM_0D = 256'h000000FFFF00000000000000000000000080007FFF8000000000000000000000;
defparam prom_inst_4.INIT_RAM_0E = 256'h0000000000000080000000FFFF80000000000000000000000000007FFFC00000;
defparam prom_inst_4.INIT_RAM_0F = 256'h000000FFFFC000000000000000000000000000FFFFC00000000001FFFF800000;
defparam prom_inst_4.INIT_RAM_10 = 256'h0100000000000020000000FFFFE00000000001FFFF8000000000000000400000;
defparam prom_inst_4.INIT_RAM_11 = 256'h000001FFFFF00000000003FFFFC000000000000000000000000001FFFFE00000;
defparam prom_inst_4.INIT_RAM_12 = 256'h000007FFFFC000000000000000000000000001FFFFE000000000000000100000;
defparam prom_inst_4.INIT_RAM_13 = 256'h0000000000000000040003FFFFF000000000000000000000000001FFFFF00000;
defparam prom_inst_4.INIT_RAM_14 = 256'h000007FFFFF000000000000000000000000003FFFFF80000000007FFFFE00000;
defparam prom_inst_4.INIT_RAM_15 = 256'h0000000000000000000007FFFFF8000000000FFFFFF000000000000000000010;
defparam prom_inst_4.INIT_RAM_16 = 256'h000007FFFFFC000000001FFFFFF000000000000000000000000007FFFFF80000;
defparam prom_inst_4.INIT_RAM_17 = 256'h00001FFFFFF80000000000000000000000000FFFFFFC00000800000000000004;
defparam prom_inst_4.INIT_RAM_18 = 256'h000000000000000000000FFFFFFC0000000000000002000000000FFFFFFE0000;
defparam prom_inst_4.INIT_RAM_19 = 256'h20001FFFFFFE0000000020000000000000000FFFFFFE000000003FFFFFF80000;
defparam prom_inst_4.INIT_RAM_1A = 256'h000000000000000000001FFFFFFF000000003FFFFFFC00000000000000000000;
defparam prom_inst_4.INIT_RAM_1B = 256'h00003FFFFFFF000000007FFFFFFE0000000000000000000200003FFFFFFE0000;
defparam prom_inst_4.INIT_RAM_1C = 256'h0000FFFFFFFE0000000000000000000000003FFFFFFF00000000000000000000;
defparam prom_inst_4.INIT_RAM_1D = 256'h000000000000000000007FFFFFFF8000400000000000000080003FFFFFFF8000;
defparam prom_inst_4.INIT_RAM_1E = 256'h00007FFFFFFF8000000000000000400000007FFFFFFF80000000FFFFFFFF0000;
defparam prom_inst_4.INIT_RAM_1F = 256'h000100000000000000007FFFFFFFC0000001FFFFFFFF00000000000000000000;
defparam prom_inst_4.INIT_RAM_20 = 256'h0000FFFFFFFFE0000001FFFFFFFF800000000000000000000000FFFFFFFFC000;
defparam prom_inst_4.INIT_RAM_21 = 256'h0003FFFFFFFFC00000000000000000000001FFFFFFFFE0000000000000000000;
defparam prom_inst_4.INIT_RAM_22 = 256'h00000000000000000001FFFFFFFFE00000000000000000000001FFFFFFFFE000;
defparam prom_inst_4.INIT_RAM_23 = 256'h0003FFFFFFFFF00000000000000000000001FFFFFFFFF0000007FFFFFFFFC000;
defparam prom_inst_4.INIT_RAM_24 = 256'h00000000000008000003FFFFFFFFF0000007FFFFFFFFE0000000000000000000;
defparam prom_inst_4.INIT_RAM_25 = 256'h0003FFFFFFFFF800000FFFFFFFFFE00000000000000000000007FFFFFFFFF000;
defparam prom_inst_4.INIT_RAM_26 = 256'h001FFFFFFFFFF00000000000000000000007FFFFFFFFF8000008000000000000;
defparam prom_inst_4.INIT_RAM_27 = 256'h0000000000000000000FFFFFFFFFFC0000000000000000000007FFFFFFFFFC00;
defparam prom_inst_4.INIT_RAM_28 = 256'h001FFFFFFFFFFC000000000000000000000FFFFFFFFFFC00001FFFFFFFFFF800;
defparam prom_inst_4.INIT_RAM_29 = 256'h0000000000000000000FFFFFFFFFFE00003FFFFFFFFFF8000000000000000000;
defparam prom_inst_4.INIT_RAM_2A = 256'h001FFFFFFFFFFC00003FFFFFFFFFFC000000000000000000001FFFFFFFFFFE00;
defparam prom_inst_4.INIT_RAM_2B = 256'h003FFFFFFFFFFC000000000000000000003FFFFFFFFFFE000000000000000100;
defparam prom_inst_4.INIT_RAM_2C = 256'h0000000000000000003FFFFFFFFFFF000000000000000000001FFFFFFFFFFC00;
defparam prom_inst_4.INIT_RAM_2D = 256'h007FFFFFFFFFFF800000000000000080003FFFFFFFFFF800003FFFFFFFFFFE00;
defparam prom_inst_4.INIT_RAM_2E = 256'h0080000000000000003FFFFFFFFFF000001FFFFFFFFFFE000000000000000000;
defparam prom_inst_4.INIT_RAM_2F = 256'h007FFFFFFFFFF000000FFFFFFFFFFF000000000000000000007FFFFFFFFFFF80;
defparam prom_inst_4.INIT_RAM_30 = 256'h000FFFFFFFFFFF80008000000000000000FFFFFFFFFFFFC00000000000000000;
defparam prom_inst_4.INIT_RAM_31 = 256'h000000000000010001FFFFFFFFFFFFC0000000000000000000FFFFFFFFFFE000;
defparam prom_inst_4.INIT_RAM_32 = 256'h01FFFFFFFFFFFFE0000000000000000000FFFFFFFFFFE0000007FFFFFFFFFF80;
defparam prom_inst_4.INIT_RAM_33 = 256'h000000000000000001FFFFFFFFFFC0000007FFFFFFFFFFC00000000000000000;
defparam prom_inst_4.INIT_RAM_34 = 256'h01FFFFFFFFFF80000003FFFFFFFFFFC0000000000000000003FFFFFFFFFFFFF0;
defparam prom_inst_4.INIT_RAM_35 = 256'h0001FFFFFFFFFFE0000000000000000003FFFFFFFFFFFFF00000000000000000;
defparam prom_inst_4.INIT_RAM_36 = 256'h001000000000000007FFFFFFFFFFFFF8000000000000000003FFFFFFFFFF8000;
defparam prom_inst_4.INIT_RAM_37 = 256'h0FFFFFFFFFFFFFF8000000000000000007FFFFFFFFFF00000001FFFFFFFFFFF0;
defparam prom_inst_4.INIT_RAM_38 = 256'h000000000000000007FFFFFFFFFF00000000FFFFFFFFFFF00000000000000800;
defparam prom_inst_4.INIT_RAM_39 = 256'h0FFFFFFFFFFE00000000FFFFFFFFFFF800000000000000000FFFFFFFFFFFFFFC;
defparam prom_inst_4.INIT_RAM_3A = 256'h00007FFFFFFFFFF800000000000000001FFFFFFFFFFFFFFE0000000000000000;
defparam prom_inst_4.INIT_RAM_3B = 256'h00000000000000001FFFFFFFFFFFFFFE00000000000000000FFFFFFFFFFC0000;
defparam prom_inst_4.INIT_RAM_3C = 256'h3FFFFFFFFFFFFFFF00000000000000001FFFFFFFFFFC000000003FFFFFFFFFFC;
defparam prom_inst_4.INIT_RAM_3D = 256'h00000000000000003FFFFFFFFFF8000000003FFFFFFFFFFE0002000000000000;
defparam prom_inst_4.INIT_RAM_3E = 256'h3FFFFFFFFFF8000000001FFFFFFFFFFE00000000000040007FFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_3F = 256'h00001FFFFFFFFFFF00000000000000007FFFFFFFFFFFFFFF8000000000000000;

pROM prom_inst_5 (
    .DO({prom_inst_5_dout_w[30:0],prom_inst_5_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_11),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_5.READ_MODE = 1'b0;
defparam prom_inst_5.BIT_WIDTH = 1;
defparam prom_inst_5.RESET_MODE = "SYNC";
defparam prom_inst_5.INIT_RAM_00 = 256'h0000000000000000FFFFFFFFFFFFFFFFC0000000000000007FFFFFFFFFF00000;
defparam prom_inst_5.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFC0000000000000007FFFFFFFFFE0000000000FFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_02 = 256'hE000000000000000FFFFFFFFFFE00000000007FFFFFFFFFF8000000000000000;
defparam prom_inst_5.INIT_RAM_03 = 256'hFFFFFFFFFFC00000000007FFFFFFFFFFC000400000000001FFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_04 = 256'h000003FFFFFFFFFFC000000000020003FFFFFFFFFFFFFFFFE000000000000001;
defparam prom_inst_5.INIT_RAM_05 = 256'hE000000000000003FFFFFFFFFFFFFFFFF000000000000001FFFFFFFFFFC00000;
defparam prom_inst_5.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFF800000000000003FFFFFFFFFF800000000003FFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_07 = 256'hF800000000000003FFFFFFFFFF000000000001FFFFFFFFFFE000000000000007;
defparam prom_inst_5.INIT_RAM_08 = 256'hFFFFFFFFFF000000000000FFFFFFFFFFF000000000000007FFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_09 = 256'h000000FFFFFFFFFFF80008000000000FFFFFFFFFFFFFFFFFFC00000000000007;
defparam prom_inst_5.INIT_RAM_0A = 256'hF80000000010001FFFFFFFFFFFFFFFFFFC0000000000000FFFFFFFFFFE000000;
defparam prom_inst_5.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFE0000000000000FFFFFFFFFFE0000000000007FFFFFFFFF;
defparam prom_inst_5.INIT_RAM_0C = 256'hFF0000000000001FFFFFFFFFFC0000000000007FFFFFFFFFFC0000000000001F;
defparam prom_inst_5.INIT_RAM_0D = 256'hFFFFFFFFF80000000000003FFFFFFFFFFC0000000000003FFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_0E = 256'h0000001FFFFFFFFFFE0000000040003FFFFFFFFFFFFFFFFFFF0000000000001F;
defparam prom_inst_5.INIT_RAM_0F = 256'hFF0001000000007FFFFFFFFFFFFFFFFFFF8000000000003FFFFFFFFFF8000000;
defparam prom_inst_5.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFF8000000000007FFFFFFFFFF00000000000001FFFFFFFFF;
defparam prom_inst_5.INIT_RAM_11 = 256'hFFC000000000007FFFFFFFFFF00000000000000FFFFFFFFFFF000000000000FF;
defparam prom_inst_5.INIT_RAM_12 = 256'hFFFFFFFFE00000000000000FFFFFFFFFFF800080000000FFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_13 = 256'h00000007FFFFFFFFFF800000000001FFFFFFFFFFFFFFFFFFFFC00000000000FF;
defparam prom_inst_5.INIT_RAM_14 = 256'hFFC00000000001FFFFFFFFFFFFFFFFFFFFE00020000001FFFFFFFFFFE0000000;
defparam prom_inst_5.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFF00000000001FFFFFFFFFFC000000000000007FFFFFFFF;
defparam prom_inst_5.INIT_RAM_16 = 256'hFFF00000000003FFFFFFFFFF8000000000000003FFFFFFFFFFE00000000003FF;
defparam prom_inst_5.INIT_RAM_17 = 256'hFFFFFFFF8000000000000001FFFFFFFFFFE00000000007FFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_18 = 256'h00000001FFFFFFFFFFF00010000007FFFFFFFFFFFFFFFFFFFFF80000000003FF;
defparam prom_inst_5.INIT_RAM_19 = 256'hFFF0000000000FFFFFFFFFFF7FFFFFFFFFF80000000007FFFFFFFFFF00000000;
defparam prom_inst_5.INIT_RAM_1A = 256'hFFFFFFFE3FFFFFFFFFFC000400000FFFFFFFFFFF0000000000000000FFFFFFFF;
defparam prom_inst_5.INIT_RAM_1B = 256'hFFFE000000000FFFFFFFFFFE0000000000000000FFFFFFFFFFF8000000000FFF;
defparam prom_inst_5.INIT_RAM_1C = 256'hFFFFFFFE00000000000000007FFFFFFFFFFC000000001FFFFFFFFFFE3FFFFFFF;
defparam prom_inst_5.INIT_RAM_1D = 256'h000000003FFFFFFFFFFC000000003FFFFFFFFFFC1FFFFFFFFFFE000000001FFF;
defparam prom_inst_5.INIT_RAM_1E = 256'hFFFE000200003FFFFFFFFFFC0FFFFFFFFFFF000000001FFFFFFFFFFC00000000;
defparam prom_inst_5.INIT_RAM_1F = 256'hFFFFFFF80FFFFFFFFFFF000000003FFFFFFFFFF800000000000000003FFFFFFF;
defparam prom_inst_5.INIT_RAM_20 = 256'hFFFF800000007FFFFFFFFFF800000000000000001FFFFFFFFFFE000000007FFF;
defparam prom_inst_5.INIT_RAM_21 = 256'hFFFFFFF000000000000000001FFFFFFFFFFF000000007FFFFFFFFFF007FFFFFF;
defparam prom_inst_5.INIT_RAM_22 = 256'h000000000FFFFFFFFFFF80000000FFFFFFFFFFF007FFFFFFFFFFC00000007FFF;
defparam prom_inst_5.INIT_RAM_23 = 256'hFFFF80000001FFFFFFFFFFE003FFFFFFFFFFC0000000FFFFFFFFFFE000000000;
defparam prom_inst_5.INIT_RAM_24 = 256'hFFFFFFE001FFFFFFFFFFE0000000FFFFFFFFFFE0000000000000000007FFFFFF;
defparam prom_inst_5.INIT_RAM_25 = 256'hFFFFE0000001FFFFFFFFFFC0000000000000000007FFFFFFFFFFC0000001FFFF;
defparam prom_inst_5.INIT_RAM_26 = 256'hFFFFFFC0000000000000000003FFFFFFFFFFC0000003FFFFFFFFFFC001FFFFFF;
defparam prom_inst_5.INIT_RAM_27 = 256'h0000000001FFFFFFFFFFE0000003FFFFFFFFFF8000FFFFFFFFFFF0000003FFFF;
defparam prom_inst_5.INIT_RAM_28 = 256'hFFFFF0000007FFFFFFFFFF8000FFFFFFFFFFF8000003FFFFFFFFFF8000000000;
defparam prom_inst_5.INIT_RAM_29 = 256'hFFFFFF00007FFFFFFFFFF8000007FFFFFFFFFF00000000000000000001FFFFFF;
defparam prom_inst_5.INIT_RAM_2A = 256'hFFFFFC000007FFFFFFFFFF00000000000000000000FFFFFFFFFFF000000FFFFF;
defparam prom_inst_5.INIT_RAM_2B = 256'hFFFFFE00000000000000000000FFFFFFFFFFF800000FFFFFFFFFFF00003FFFFF;
defparam prom_inst_5.INIT_RAM_2C = 256'h00000000007FFFFFFFFFF800001FFFFFFFFFFE00003FFFFFFFFFFE00000FFFFF;
defparam prom_inst_5.INIT_RAM_2D = 256'hFFFFFC00003FFFFFFFFFFC00001FFFFFFFFFFE00001FFFFFFFFFFE0000000000;
defparam prom_inst_5.INIT_RAM_2E = 256'hFFFFFC00001FFFFFFFFFFF00001FFFFFFFFFFC000000000000000000003FFFFF;
defparam prom_inst_5.INIT_RAM_2F = 256'hFFFFFF00003FFFFFFFFFF8000000000000000000003FFFFFFFFFFE00003FFFFF;
defparam prom_inst_5.INIT_RAM_30 = 256'hFFFFF8000000000000000000001FFFFFFFFFFE00007FFFFFFFFFF800000FFFFF;
defparam prom_inst_5.INIT_RAM_31 = 256'h00000000001FFFFFFFFFFF00007FFFFFFFFFF8000007FFFFFFFFFF80003FFFFF;
defparam prom_inst_5.INIT_RAM_32 = 256'hFFFFFF0000FFFFFFFFFFF0000007FFFFFFFFFFC0007FFFFFFFFFF00000000000;
defparam prom_inst_5.INIT_RAM_33 = 256'hFFFFE0000003FFFFFFFFFFC000FFFFFFFFFFF0000000000000000000000FFFFF;
defparam prom_inst_5.INIT_RAM_34 = 256'hFFFFFFE000FFFFFFFFFFE00000000000000000000007FFFFFFFFFF8001FFFFFF;
defparam prom_inst_5.INIT_RAM_35 = 256'hFFFFE00000000000000000000007FFFFFFFFFFC001FFFFFFFFFFE0000003FFFF;
defparam prom_inst_5.INIT_RAM_36 = 256'h000000000003FFFFFFFFFFC003FFFFFFFFFFC0000001FFFFFFFFFFE001FFFFFF;
defparam prom_inst_5.INIT_RAM_37 = 256'hFFFFFFE003FFFFFFFFFFC0000001FFFFFFFFFFF001FFFFFFFFFFC00000000000;
defparam prom_inst_5.INIT_RAM_38 = 256'hFFFF80000000FFFFFFFFFFF003FFFFFFFFFF800000000000000000000003FFFF;
defparam prom_inst_5.INIT_RAM_39 = 256'hFFFFFFF803FFFFFFFFFF800000000000000000000001FFFFFFFFFFE007FFFFFF;
defparam prom_inst_5.INIT_RAM_3A = 256'hFFFF000000000000000000000000FFFFFFFFFFF00FFFFFFFFFFF000000007FFF;
defparam prom_inst_5.INIT_RAM_3B = 256'h000000000000FFFFFFFFFFF00FFFFFFFFFFF000000007FFFFFFFFFFC07FFFFFF;
defparam prom_inst_5.INIT_RAM_3C = 256'hFFFFFFF81FFFFFFFFFFE000000003FFFFFFFFFFC0FFFFFFFFFFF000000000000;
defparam prom_inst_5.INIT_RAM_3D = 256'hFFFE000000001FFFFFFFFFFE0FFFFFFFFFFE0000000000000000000000007FFF;
defparam prom_inst_5.INIT_RAM_3E = 256'hFFFFFFFE1FFFFFFFFFFC0000000000000000000000007FFFFFFFFFFC1FFFFFFF;
defparam prom_inst_5.INIT_RAM_3F = 256'hFFFC0000000000000000000000003FFFFFFFFFFC3FFFFFFFFFFC000000001FFF;

pROM prom_inst_6 (
    .DO({prom_inst_6_dout_w[30:0],prom_inst_6_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_13),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_6.READ_MODE = 1'b0;
defparam prom_inst_6.BIT_WIDTH = 1;
defparam prom_inst_6.RESET_MODE = "SYNC";
defparam prom_inst_6.INIT_RAM_00 = 256'h0000000000001FFFFFFFFFFE7FFFFFFFFFF8000000000FFFFFFFFFFF1FFFFFFF;
defparam prom_inst_6.INIT_RAM_01 = 256'hFFFFFFFE7FFFFFFFFFF8000000000FFFFFFFFFFFBFFFFFFFFFF8000000000000;
defparam prom_inst_6.INIT_RAM_02 = 256'hFFF00000000007FFFFFFFFFFFFFFFFFFFFF80000000000000000000000001FFF;
defparam prom_inst_6.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFF00000000000000000000000000FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_04 = 256'hFFE00000000000000000000000000FFFFFFFFFFFFFFFFFFFFFE00000000003FF;
defparam prom_inst_6.INIT_RAM_05 = 256'h00000000000007FFFFFFFFFFFFFFFFFFFFE00000000003FFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFC00000000001FFFFFFFFFFFFFFFFFFFFE0000000000000;
defparam prom_inst_6.INIT_RAM_07 = 256'hFFC00000000001FFFFFFFFFFFFFFFFFFFFC000000000000000000000000003FF;
defparam prom_inst_6.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFC000000000000000000000000003FFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_09 = 256'hFF8000000000000000000000000001FFFFFFFFFFFFFFFFFFFF800000000000FF;
defparam prom_inst_6.INIT_RAM_0A = 256'h00000000000001FFFFFFFFFFFFFFFFFFFF0000000000007FFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFF0000000000007FFFFFFFFFFFFFFFFFFF00000000000000;
defparam prom_inst_6.INIT_RAM_0C = 256'hFE0000000000003FFFFFFFFFFFFFFFFFFF0000000000000000000000000000FF;
defparam prom_inst_6.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFE00000000000000000000000000007FFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_0E = 256'hFE00000000000000000000000000007FFFFFFFFFFFFFFFFFFE0000000000003F;
defparam prom_inst_6.INIT_RAM_0F = 256'h000000000000003FFFFFFFFFFFFFFFFFFC0000000000001FFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFF80000000000000FFFFFFFFFFFFFFFFFFC00000000000000;
defparam prom_inst_6.INIT_RAM_11 = 256'hF80000000000000FFFFFFFFFFFFFFFFFF800000000000000000000000000003F;
defparam prom_inst_6.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFF800000000000000000000000000001FFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_13 = 256'hF000000000000000000000000000000FFFFFFFFFFFFFFFFFF000000000000007;
defparam prom_inst_6.INIT_RAM_14 = 256'h000000000000000FFFFFFFFFFFFFFFFFF000000000000007FFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFE000000000000003FFFFFFFFFFFFFFFFF000000000000000;
defparam prom_inst_6.INIT_RAM_16 = 256'hC000000000000001FFFFFFFFFFFFFFFFE0000000000000000000000000000007;
defparam prom_inst_6.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFE0000000000000000000000000000007FFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_18 = 256'hC0000000000000000000000000000003FFFFFFFFFFFFFFFFC000000000000001;
defparam prom_inst_6.INIT_RAM_19 = 256'h0000000000000001FFFFFFFFFFFFFFFF8000000000000000FFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFF8000000000000000FFFFFFFFFFFFFFFF8000000000000000;
defparam prom_inst_6.INIT_RAM_1B = 256'h00000000000000007FFFFFFFFFFFFFFF80000000000000000000000000000001;
defparam prom_inst_6.INIT_RAM_1C = 256'h7FFFFFFFFFFFFFFF00000000000000000000000000000000FFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1D = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFF0000000000000000;
defparam prom_inst_6.INIT_RAM_1E = 256'h00000000000000007FFFFFFFFFFFFFFE00000000000000003FFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1F = 256'h7FFFFFFFFFFFFFFC00000000000000001FFFFFFFFFFFFFFE0000000000000000;
defparam prom_inst_6.INIT_RAM_20 = 256'h00000000000000001FFFFFFFFFFFFFFC00000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_21 = 256'h0FFFFFFFFFFFFFFC000000000000000000000000000000003FFFFFFFFFFFFFFC;
defparam prom_inst_6.INIT_RAM_22 = 256'h000000000000000000000000000000001FFFFFFFFFFFFFF80000000000000000;
defparam prom_inst_6.INIT_RAM_23 = 256'h00000000000000001FFFFFFFFFFFFFF800000000000000000FFFFFFFFFFFFFF8;
defparam prom_inst_6.INIT_RAM_24 = 256'h0FFFFFFFFFFFFFF0000000000000000007FFFFFFFFFFFFF80000000000000000;
defparam prom_inst_6.INIT_RAM_25 = 256'h000000000000000003FFFFFFFFFFFFF000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_26 = 256'h03FFFFFFFFFFFFF0000000000000000000000000000000000FFFFFFFFFFFFFE0;
defparam prom_inst_6.INIT_RAM_27 = 256'h0000000000000000000000000000000007FFFFFFFFFFFFE00000000000000000;
defparam prom_inst_6.INIT_RAM_28 = 256'h000000000000000003FFFFFFFFFFFFC0000000000000000001FFFFFFFFFFFFE0;
defparam prom_inst_6.INIT_RAM_29 = 256'h03FFFFFFFFFFFFC0000000000000000001FFFFFFFFFFFFC00000000000000000;
defparam prom_inst_6.INIT_RAM_2A = 256'h000000000000000000FFFFFFFFFFFFC000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_2B = 256'h007FFFFFFFFFFF800000000000000000000000000000000001FFFFFFFFFFFF80;
defparam prom_inst_6.INIT_RAM_2C = 256'h0000000000000000000000000000000000FFFFFFFFFFFF000000000000000000;
defparam prom_inst_6.INIT_RAM_2D = 256'h000000000000000000FFFFFFFFFFFF000000000000000000007FFFFFFFFFFF00;
defparam prom_inst_6.INIT_RAM_2E = 256'h007FFFFFFFFFFE000000000000000000003FFFFFFFFFFF000000000000000000;
defparam prom_inst_6.INIT_RAM_2F = 256'h0000000000000000003FFFFFFFFFFE0000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_30 = 256'h001FFFFFFFFFFE0000000000000000000000000000000000007FFFFFFFFFFE00;
defparam prom_inst_6.INIT_RAM_31 = 256'h00000000000000000000000000000000003FFFFFFFFFFC000000000000000000;
defparam prom_inst_6.INIT_RAM_32 = 256'h0000000000000000001FFFFFFFFFF8000000000000000000000FFFFFFFFFFC00;
defparam prom_inst_6.INIT_RAM_33 = 256'h001FFFFFFFFFF8000000000000000000000FFFFFFFFFF8000000000000000000;
defparam prom_inst_6.INIT_RAM_34 = 256'h00000000000000000007FFFFFFFFF80000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_35 = 256'h0007FFFFFFFFF00000000000000000000000000000000000000FFFFFFFFFF000;
defparam prom_inst_6.INIT_RAM_36 = 256'h00000000000000000000000000000000000FFFFFFFFFF0000000000000000000;
defparam prom_inst_6.INIT_RAM_37 = 256'h00000000000000000007FFFFFFFFE00000000000000000000003FFFFFFFFF000;
defparam prom_inst_6.INIT_RAM_38 = 256'h0003FFFFFFFFC00000000000000000000001FFFFFFFFE0000000000000000000;
defparam prom_inst_6.INIT_RAM_39 = 256'h00000000000000000001FFFFFFFFC00000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_3A = 256'h0000FFFFFFFFC000000000000000000000000000000000000003FFFFFFFFC000;
defparam prom_inst_6.INIT_RAM_3B = 256'h000000000000000000000000000000000001FFFFFFFF80000000000000000000;
defparam prom_inst_6.INIT_RAM_3C = 256'h00000000000000000001FFFFFFFF800000000000000000000000FFFFFFFF8000;
defparam prom_inst_6.INIT_RAM_3D = 256'h0000FFFFFFFF0000000000000000000000007FFFFFFF80000000000000000000;
defparam prom_inst_6.INIT_RAM_3E = 256'h000000000000000000003FFFFFFF000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_3F = 256'h00003FFFFFFF00000000000000000000000000000000000000007FFFFFFE0000;

pROM prom_inst_7 (
    .DO({prom_inst_7_dout_w[30:0],prom_inst_7_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_15),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_7.READ_MODE = 1'b0;
defparam prom_inst_7.BIT_WIDTH = 1;
defparam prom_inst_7.RESET_MODE = "SYNC";
defparam prom_inst_7.INIT_RAM_00 = 256'h0000000000000000000000000000000000007FFFFFFE00000000000000000000;
defparam prom_inst_7.INIT_RAM_01 = 256'h000000000000000000003FFFFFFC0000000000000000000000001FFFFFFE0000;
defparam prom_inst_7.INIT_RAM_02 = 256'h00003FFFFFFC0000000000000000000000001FFFFFFC00000000000000000000;
defparam prom_inst_7.INIT_RAM_03 = 256'h000000000000000000000FFFFFFC000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_04 = 256'h00000FFFFFF800000000000000000000000000000000000000001FFFFFF80000;
defparam prom_inst_7.INIT_RAM_05 = 256'h0000000000000000000000000000000000000FFFFFF000000000000000000000;
defparam prom_inst_7.INIT_RAM_06 = 256'h000000000000000000000FFFFFF000000000000000000000000007FFFFF80000;
defparam prom_inst_7.INIT_RAM_07 = 256'h000007FFFFE000000000000000000000000003FFFFF000000000000000000000;
defparam prom_inst_7.INIT_RAM_08 = 256'h0000000000000000000001FFFFE0000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_09 = 256'h000001FFFFE0000000000000000000000000000000000000000007FFFFC00000;
defparam prom_inst_7.INIT_RAM_0A = 256'h00000000000000000000000000000000000003FFFFC000000000000000000000;
defparam prom_inst_7.INIT_RAM_0B = 256'h0000000000000000000001FFFF8000000000000000000000000000FFFFC00000;
defparam prom_inst_7.INIT_RAM_0C = 256'h000001FFFF8000000000000000000000000000FFFFC000000000000000000000;
defparam prom_inst_7.INIT_RAM_0D = 256'h00000000000000000000007FFF80000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_0E = 256'h0000003FFF00000000000000000000000000000000000000000000FFFF000000;
defparam prom_inst_7.INIT_RAM_0F = 256'h00000000000000000000000000000000000000FFFE0000000000000000000000;
defparam prom_inst_7.INIT_RAM_10 = 256'h00000000000000000000007FFE00000000000000000000000000003FFF000000;
defparam prom_inst_7.INIT_RAM_11 = 256'h0000003FFC00000000000000000000000000001FFE0000000000000000000000;
defparam prom_inst_7.INIT_RAM_12 = 256'h00000000000000000000001FFE00000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_13 = 256'h0000000FFC000000000000000000000000000000000000000000003FFC000000;
defparam prom_inst_7.INIT_RAM_14 = 256'h000000000000000000000000000000000000001FF80000000000000000000000;
defparam prom_inst_7.INIT_RAM_15 = 256'h00000000000000000000001FF0000000000000000000000000000007F8000000;
defparam prom_inst_7.INIT_RAM_16 = 256'h0000000FF0000000000000000000000000000007F80000000000000000000000;
defparam prom_inst_7.INIT_RAM_17 = 256'h000000000000000000000003F000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_18 = 256'h00000003F00000000000000000000000000000000000000000000007E0000000;
defparam prom_inst_7.INIT_RAM_19 = 256'h0000000000000000000000000000000000000007E00000000000000000000000;
defparam prom_inst_7.INIT_RAM_1A = 256'h000000000000000000000003C0000000000000000000000000000001E0000000;
defparam prom_inst_7.INIT_RAM_1B = 256'h0000000380000000000000000000000000000001E00000000000000000000000;
defparam prom_inst_7.INIT_RAM_1C = 256'h000000000000000000000000C000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000180000000;
defparam prom_inst_7.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_8 (
    .DO({prom_inst_8_dout_w[30:0],prom_inst_8_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_8.READ_MODE = 1'b0;
defparam prom_inst_8.BIT_WIDTH = 1;
defparam prom_inst_8.RESET_MODE = "SYNC";
defparam prom_inst_8.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_9 (
    .DO({prom_inst_9_dout_w[30:0],prom_inst_9_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_3),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_9.READ_MODE = 1'b0;
defparam prom_inst_9.BIT_WIDTH = 1;
defparam prom_inst_9.RESET_MODE = "SYNC";
defparam prom_inst_9.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_37 = 256'h0000000000000000000000008000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_38 = 256'h0000000180000000000000000000000000000000C00000000000000000000000;
defparam prom_inst_9.INIT_RAM_39 = 256'h000000000000000000000001C000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_3A = 256'h00000001E00000000000000000000000000000000000000000000001C0000000;
defparam prom_inst_9.INIT_RAM_3B = 256'h0000000000000000000000000000000000000003C00000000000000000000000;
defparam prom_inst_9.INIT_RAM_3C = 256'h000000000000000000000007E0000000000000000000000000000003F0000000;
defparam prom_inst_9.INIT_RAM_3D = 256'h00000007F0000000000000000000000000000003F00000000000000000000000;
defparam prom_inst_9.INIT_RAM_3E = 256'h000000000000000000000007F800000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_3F = 256'h0000000FF8000000000000000000000000000000000000000000000FF0000000;

pROM prom_inst_10 (
    .DO({prom_inst_10_dout_w[30:0],prom_inst_10_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_5),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_10.READ_MODE = 1'b0;
defparam prom_inst_10.BIT_WIDTH = 1;
defparam prom_inst_10.RESET_MODE = "SYNC";
defparam prom_inst_10.INIT_RAM_00 = 256'h000000000000000000000000000000000000000FF80000000000000000000000;
defparam prom_inst_10.INIT_RAM_01 = 256'h00000000000000000000001FF800000000000000000000000000000FFC000000;
defparam prom_inst_10.INIT_RAM_02 = 256'h0000003FFC00000000000000000000000000001FFE0000000000000000000000;
defparam prom_inst_10.INIT_RAM_03 = 256'h00000000000000000000001FFE00000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_04 = 256'h0000003FFF000000000000000000000000000000000000000000003FFE000000;
defparam prom_inst_10.INIT_RAM_05 = 256'h000000000000000000000000000000000000007FFE0000000000000000000000;
defparam prom_inst_10.INIT_RAM_06 = 256'h00000000000000000000007FFF00000000000000000000000000007FFF000000;
defparam prom_inst_10.INIT_RAM_07 = 256'h000000FFFF00000000000000000000000000007FFF8000000000000000000000;
defparam prom_inst_10.INIT_RAM_08 = 256'h0000000000000000000000FFFFC0000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_09 = 256'h000000FFFFC0000000000000000000000000000000000000000001FFFF800000;
defparam prom_inst_10.INIT_RAM_0A = 256'h00000000000000000000000000000000000001FFFFC000000000000000000000;
defparam prom_inst_10.INIT_RAM_0B = 256'h0000000000000000000003FFFFC000000000000000000000000001FFFFE00000;
defparam prom_inst_10.INIT_RAM_0C = 256'h000003FFFFE000000000000000000000000003FFFFE000000000000000000000;
defparam prom_inst_10.INIT_RAM_0D = 256'h0000000000000000000003FFFFF0000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_0E = 256'h000007FFFFF8000000000000000000000000000000000000000007FFFFF00000;
defparam prom_inst_10.INIT_RAM_0F = 256'h0000000000000000000000000000000000000FFFFFF000000000000000000000;
defparam prom_inst_10.INIT_RAM_10 = 256'h000000000000000000000FFFFFF80000000000000000000000000FFFFFF80000;
defparam prom_inst_10.INIT_RAM_11 = 256'h00001FFFFFF80000000000000000000000000FFFFFFC00000000000000000000;
defparam prom_inst_10.INIT_RAM_12 = 256'h000000000000000000001FFFFFFC000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_13 = 256'h00001FFFFFFE00000000000000000000000000000000000000001FFFFFFC0000;
defparam prom_inst_10.INIT_RAM_14 = 256'h0000000000000000000000000000000000003FFFFFFE00000000000000000000;
defparam prom_inst_10.INIT_RAM_15 = 256'h000000000000000000007FFFFFFE0000000000000000000000003FFFFFFF0000;
defparam prom_inst_10.INIT_RAM_16 = 256'h00007FFFFFFF0000000000000000000000007FFFFFFF00000000000000000000;
defparam prom_inst_10.INIT_RAM_17 = 256'h000000000000000000007FFFFFFF800000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_18 = 256'h0000FFFFFFFF8000000000000000000000000000000000000000FFFFFFFF0000;
defparam prom_inst_10.INIT_RAM_19 = 256'h000000000000000000000000000000000000FFFFFFFF80000000000000000000;
defparam prom_inst_10.INIT_RAM_1A = 256'h00000000000000000001FFFFFFFF800000000000000000000000FFFFFFFFC000;
defparam prom_inst_10.INIT_RAM_1B = 256'h0001FFFFFFFFC00000000000000000000001FFFFFFFFC0000000000000000000;
defparam prom_inst_10.INIT_RAM_1C = 256'h00000000000000000001FFFFFFFFE00000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_1D = 256'h0003FFFFFFFFF000000000000000000000000000000000000003FFFFFFFFE000;
defparam prom_inst_10.INIT_RAM_1E = 256'h000000000000000000000000000000000007FFFFFFFFE0000000000000000000;
defparam prom_inst_10.INIT_RAM_1F = 256'h00000000000000000007FFFFFFFFF00000000000000000000007FFFFFFFFF000;
defparam prom_inst_10.INIT_RAM_20 = 256'h000FFFFFFFFFF00000000000000000000007FFFFFFFFF8000000000000000000;
defparam prom_inst_10.INIT_RAM_21 = 256'h0000000000000000000FFFFFFFFFF80000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_22 = 256'h000FFFFFFFFFFC0000000000000000000000000000000000000FFFFFFFFFF800;
defparam prom_inst_10.INIT_RAM_23 = 256'h00000000000000000000000000000000001FFFFFFFFFFC000000000000000000;
defparam prom_inst_10.INIT_RAM_24 = 256'h0000000000000000003FFFFFFFFFFC000000000000000000001FFFFFFFFFFE00;
defparam prom_inst_10.INIT_RAM_25 = 256'h003FFFFFFFFFFE000000000000000000003FFFFFFFFFFE000000000000000000;
defparam prom_inst_10.INIT_RAM_26 = 256'h0000000000000000003FFFFFFFFFFF0000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_27 = 256'h007FFFFFFFFFFF0000000000000000000000000000000000007FFFFFFFFFFE00;
defparam prom_inst_10.INIT_RAM_28 = 256'h00000000000000000000000000000000007FFFFFFFFFFF000000000000000000;
defparam prom_inst_10.INIT_RAM_29 = 256'h000000000000000000FFFFFFFFFFFF800000000000000000007FFFFFFFFFFF80;
defparam prom_inst_10.INIT_RAM_2A = 256'h007FFFFFFFFFFF000000000000000000007FFFFFFFFFFF800000000000000000;
defparam prom_inst_10.INIT_RAM_2B = 256'h0000000000000000003FFFFFFFFFFF0000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_2C = 256'h003FFFFFFFFFFE0000000000000000000000000000000000007FFFFFFFFFFE00;
defparam prom_inst_10.INIT_RAM_2D = 256'h00000000000000000000000000000000003FFFFFFFFFFE000000000000000000;
defparam prom_inst_10.INIT_RAM_2E = 256'h0000000000000000003FFFFFFFFFFC000000000000000000001FFFFFFFFFFE00;
defparam prom_inst_10.INIT_RAM_2F = 256'h001FFFFFFFFFFC000000000000000000001FFFFFFFFFFC000000000000000000;
defparam prom_inst_10.INIT_RAM_30 = 256'h0000000000000000000FFFFFFFFFFC0000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_31 = 256'h0007FFFFFFFFF80000000000000000000000000000000000000FFFFFFFFFF800;
defparam prom_inst_10.INIT_RAM_32 = 256'h00000000000000000000000000000000000FFFFFFFFFF0000000000000000000;
defparam prom_inst_10.INIT_RAM_33 = 256'h00000000000000000007FFFFFFFFF00000000000000000000007FFFFFFFFF000;
defparam prom_inst_10.INIT_RAM_34 = 256'h0007FFFFFFFFE00000000000000000000003FFFFFFFFF0000000000000000000;
defparam prom_inst_10.INIT_RAM_35 = 256'h00000000000000000003FFFFFFFFE00000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_36 = 256'h0001FFFFFFFFE000000000000000000000000000000000000003FFFFFFFFE000;
defparam prom_inst_10.INIT_RAM_37 = 256'h000000000000000000000000000000000001FFFFFFFFC0000000000000000000;
defparam prom_inst_10.INIT_RAM_38 = 256'h00000000000000000001FFFFFFFF800000000000000000000000FFFFFFFFC000;
defparam prom_inst_10.INIT_RAM_39 = 256'h8000FFFFFFFF800080000000000000004000FFFFFFFF80000000000000000000;
defparam prom_inst_10.INIT_RAM_3A = 256'h8000000000000000C0007FFFFFFF8000C0000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_3B = 256'hE0007FFFFFFF0001C00000000000000000000000000000018000FFFFFFFF0001;
defparam prom_inst_10.INIT_RAM_3C = 256'hE0000000000000000000000000000001C0007FFFFFFF0001C000000000000000;
defparam prom_inst_10.INIT_RAM_3D = 256'h0000000000000003C0007FFFFFFE0003C000000000000001E0003FFFFFFF0001;
defparam prom_inst_10.INIT_RAM_3E = 256'hE0003FFFFFFE0003E000000000000003F0003FFFFFFE0003F000000000000000;
defparam prom_inst_10.INIT_RAM_3F = 256'hF000000000000003F0001FFFFFFE0003F0000000000000000000000000000003;

pROM prom_inst_11 (
    .DO({prom_inst_11_dout_w[30:0],prom_inst_11_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_7),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_11.READ_MODE = 1'b0;
defparam prom_inst_11.BIT_WIDTH = 1;
defparam prom_inst_11.RESET_MODE = "SYNC";
defparam prom_inst_11.INIT_RAM_00 = 256'hF8000FFFFFFC0007F8000000000000000000000000000007F0001FFFFFFC0007;
defparam prom_inst_11.INIT_RAM_01 = 256'hF800000000000000000000000000000FF0001FFFFFF8000FF000000000000007;
defparam prom_inst_11.INIT_RAM_02 = 256'h000000000000000FF8000FFFFFF8000FF800000000000007FC000FFFFFF8000F;
defparam prom_inst_11.INIT_RAM_03 = 256'hF8000FFFFFF0001FF80000000000000FFC0007FFFFF8000FFC00000000000000;
defparam prom_inst_11.INIT_RAM_04 = 256'hFC0000000000001FFE0003FFFFF0001FFE00000000000000000000000000001F;
defparam prom_inst_11.INIT_RAM_05 = 256'hFE0003FFFFF0001FFE00000000000000000000000000001FFC0007FFFFF0001F;
defparam prom_inst_11.INIT_RAM_06 = 256'hFF00000000000000000000000000003FFE0003FFFFE0003FFE0000000000001F;
defparam prom_inst_11.INIT_RAM_07 = 256'h000000000000007FFE0003FFFFC0007FFE0000000000003FFF0001FFFFE0003F;
defparam prom_inst_11.INIT_RAM_08 = 256'hFF0001FFFFC0007FFF0000000000003FFF8000FFFFC0007FFF00000000000000;
defparam prom_inst_11.INIT_RAM_09 = 256'hFF0000000000007FFF8000FFFFC0007FFF80000000000000000000000000007F;
defparam prom_inst_11.INIT_RAM_0A = 256'hFFC0007FFF8000FFFFC000000000000000000000000000FFFF8001FFFF8000FF;
defparam prom_inst_11.INIT_RAM_0B = 256'hFFC000000000000000000000000000FFFF8000FFFF0000FFFF800000000000FF;
defparam prom_inst_11.INIT_RAM_0C = 256'h00000000000001FFFFC0007FFF0001FFFFC00000000000FFFFC0007FFF0001FF;
defparam prom_inst_11.INIT_RAM_0D = 256'hFFC0007FFE0003FFFFC00000000001FFFFE0003FFF0001FFFFE0000000000000;
defparam prom_inst_11.INIT_RAM_0E = 256'hFFE00000000001FFFFF0001FFE0003FFFFE000000000000000000000000003FF;
defparam prom_inst_11.INIT_RAM_0F = 256'hFFF0001FFE0003FFFFF000000000000000000000000003FFFFE0003FFE0003FF;
defparam prom_inst_11.INIT_RAM_10 = 256'hFFF800000000000000000000000007FFFFF0003FFC0007FFFFE00000000003FF;
defparam prom_inst_11.INIT_RAM_11 = 256'h00000000000007FFFFF0001FF80007FFFFF00000000007FFFFF8000FFC0007FF;
defparam prom_inst_11.INIT_RAM_12 = 256'hFFF8000FF8000FFFFFF80000000007FFFFF8000FF8000FFFFFF8000000000000;
defparam prom_inst_11.INIT_RAM_13 = 256'hFFF8000000000FFFFFFC0007F8000FFFFFFC0000000000000000000000000FFF;
defparam prom_inst_11.INIT_RAM_14 = 256'hFFFE0003F0001FFFFFFC0000000000000000000000001FFFFFF8000FF0001FFF;
defparam prom_inst_11.INIT_RAM_15 = 256'hFFFE0000000000000000000000001FFFFFFC0007F0001FFFFFFC000000000FFF;
defparam prom_inst_11.INIT_RAM_16 = 256'h0000000000003FFFFFFE0007E0003FFFFFFE000000001FFFFFFE0003F0001FFF;
defparam prom_inst_11.INIT_RAM_17 = 256'hFFFE0003C0003FFFFFFE000000003FFFFFFF0001E0003FFFFFFF000000000000;
defparam prom_inst_11.INIT_RAM_18 = 256'hFFFF000000003FFFFFFF0001C0007FFFFFFF0000000000000000000000003FFF;
defparam prom_inst_11.INIT_RAM_19 = 256'hFFFF8000C0007FFFFFFF8000000000000000000000007FFFFFFF0001C0007FFF;
defparam prom_inst_11.INIT_RAM_1A = 256'hFFFF800000000000000000000000FFFFFFFF00018000FFFFFFFF000000007FFF;
defparam prom_inst_11.INIT_RAM_1B = 256'h000000000000FFFFFFFF80008000FFFFFFFF80000000FFFFFFFFC0000000FFFF;
defparam prom_inst_11.INIT_RAM_1C = 256'hFFFFC0000001FFFFFFFFC0000000FFFFFFFFC0000000FFFFFFFFC00000000000;
defparam prom_inst_11.INIT_RAM_1D = 256'hFFFFC0000001FFFFFFFFE0000001FFFFFFFFE00000000000000000000001FFFF;
defparam prom_inst_11.INIT_RAM_1E = 256'hFFFFE0000003FFFFFFFFE00000000000000000000001FFFFFFFFC0000001FFFF;
defparam prom_inst_11.INIT_RAM_1F = 256'hFFFFF00000000000000000000003FFFFFFFFE0000003FFFFFFFFE0000001FFFF;
defparam prom_inst_11.INIT_RAM_20 = 256'h000000000007FFFFFFFFE0000007FFFFFFFFE0000003FFFFFFFFF0000003FFFF;
defparam prom_inst_11.INIT_RAM_21 = 256'hFFFFF0000007FFFFFFFFF0000007FFFFFFFFF0000007FFFFFFFFF00000000000;
defparam prom_inst_11.INIT_RAM_22 = 256'hFFFFF0000007FFFFFFFFF8000007FFFFFFFFF80000000000000000000007FFFF;
defparam prom_inst_11.INIT_RAM_23 = 256'hFFFFFC00000FFFFFFFFFFC000000000000000000000FFFFFFFFFF800000FFFFF;
defparam prom_inst_11.INIT_RAM_24 = 256'hFFFFFC000000000000000000000FFFFFFFFFF800000FFFFFFFFFF800000FFFFF;
defparam prom_inst_11.INIT_RAM_25 = 256'h00000000001FFFFFFFFFFC00001FFFFFFFFFFC00000FFFFFFFFFFC00000FFFFF;
defparam prom_inst_11.INIT_RAM_26 = 256'hFFFFFC00003FFFFFFFFFFC00001FFFFFFFFFFE00001FFFFFFFFFFE0000000000;
defparam prom_inst_11.INIT_RAM_27 = 256'hFFFFFE00003FFFFFFFFFFF00003FFFFFFFFFFE000000000000000000001FFFFF;
defparam prom_inst_11.INIT_RAM_28 = 256'hFFFFFF00003FFFFFFFFFFF000000000000000000003FFFFFFFFFFE00003FFFFF;
defparam prom_inst_11.INIT_RAM_29 = 256'hFFFFFF800000000000000000007FFFFFFFFFFF00007FFFFFFFFFFE00003FFFFF;
defparam prom_inst_11.INIT_RAM_2A = 256'h00000000007FFFFFFFFFFF0000FFFFFFFFFFFF00007FFFFFFFFFFF80007FFFFF;
defparam prom_inst_11.INIT_RAM_2B = 256'hFFFFFF8000FFFFFFFFFFFF80007FFFFFFFFFFF80007FFFFFFFFFFF8000000000;
defparam prom_inst_11.INIT_RAM_2C = 256'hFFFFFF00007FFFFFFFFFFF80007FFFFFFFFFFF80000000000000000000FFFFFF;
defparam prom_inst_11.INIT_RAM_2D = 256'hFFFFFF00003FFFFFFFFFFF000000000000000000007FFFFFFFFFFF0000FFFFFF;
defparam prom_inst_11.INIT_RAM_2E = 256'hFFFFFE000000000000000000007FFFFFFFFFFF00007FFFFFFFFFFF00003FFFFF;
defparam prom_inst_11.INIT_RAM_2F = 256'h00000000003FFFFFFFFFFE00003FFFFFFFFFFE00003FFFFFFFFFFF00003FFFFF;
defparam prom_inst_11.INIT_RAM_30 = 256'hFFFFFC00003FFFFFFFFFFC00001FFFFFFFFFFE00001FFFFFFFFFFE0000000000;
defparam prom_inst_11.INIT_RAM_31 = 256'hFFFFFC00000FFFFFFFFFFE00001FFFFFFFFFFC000000000000000000003FFFFF;
defparam prom_inst_11.INIT_RAM_32 = 256'hFFFFFC00000FFFFFFFFFFC000000000000000000001FFFFFFFFFFC00001FFFFF;
defparam prom_inst_11.INIT_RAM_33 = 256'hFFFFF8000000000000000000000FFFFFFFFFF800000FFFFFFFFFF800000FFFFF;
defparam prom_inst_11.INIT_RAM_34 = 256'h00000000000FFFFFFFFFF800000FFFFFFFFFF8000007FFFFFFFFF8000007FFFF;
defparam prom_inst_11.INIT_RAM_35 = 256'hFFFFF0000007FFFFFFFFF0000007FFFFFFFFF8000007FFFFFFFFF00000000000;
defparam prom_inst_11.INIT_RAM_36 = 256'hFFFFE0000003FFFFFFFFF0000003FFFFFFFFF00000000000000000000007FFFF;
defparam prom_inst_11.INIT_RAM_37 = 256'hFFFFE0000003FFFFFFFFE00000000000000000000007FFFFFFFFE0000007FFFF;
defparam prom_inst_11.INIT_RAM_38 = 256'hFFFFE00000000000000000000003FFFFFFFFE0000003FFFFFFFFE0000001FFFF;
defparam prom_inst_11.INIT_RAM_39 = 256'h000000000001FFFFFFFFC0000001FFFFFFFFC0000001FFFFFFFFE0000001FFFF;
defparam prom_inst_11.INIT_RAM_3A = 256'hFFFFC0000001FFFFFFFFC0000000FFFFFFFFC0000000FFFFFFFFC00000000000;
defparam prom_inst_11.INIT_RAM_3B = 256'hFFFF80000000FFFFFFFFC0000000FFFFFFFF800000000000000000000001FFFF;
defparam prom_inst_11.INIT_RAM_3C = 256'hFFFF800080007FFFFFFF800000000000000000000000FFFFFFFF80000000FFFF;
defparam prom_inst_11.INIT_RAM_3D = 256'hFFFF000040000000000000000000FFFFFFFF00008000FFFFFFFF000000007FFF;
defparam prom_inst_11.INIT_RAM_3E = 256'h0000000180007FFFFFFF000180007FFFFFFF0000C0003FFFFFFF0000C0007FFF;
defparam prom_inst_11.INIT_RAM_3F = 256'hFFFE0001C0003FFFFFFE0000C0003FFFFFFF0001E0003FFFFFFF0000E0000000;

pROM prom_inst_12 (
    .DO({prom_inst_12_dout_w[30:0],prom_inst_12_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_9),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_12.READ_MODE = 1'b0;
defparam prom_inst_12.BIT_WIDTH = 1;
defparam prom_inst_12.RESET_MODE = "SYNC";
defparam prom_inst_12.INIT_RAM_00 = 256'hFFFE0001E0001FFFFFFE0001E0001FFFFFFE0000E00000000000000380003FFF;
defparam prom_inst_12.INIT_RAM_01 = 256'hFFFE0003F0001FFFFFFC0001F000000000000003C0003FFFFFFE0003C0003FFF;
defparam prom_inst_12.INIT_RAM_02 = 256'hFFFC0001F000000000000007C0001FFFFFFC0007E0001FFFFFFC0003F0000FFF;
defparam prom_inst_12.INIT_RAM_03 = 256'h00000007E0001FFFFFF80007F0001FFFFFF80003F0000FFFFFFC0007F0000FFF;
defparam prom_inst_12.INIT_RAM_04 = 256'hFFF8000FF0000FFFFFF00007F80007FFFFF80007F8000FFFFFF80003F8000000;
defparam prom_inst_12.INIT_RAM_05 = 256'hFFF00007F80007FFFFF8000FFC0007FFFFF80007FC0000000000000FF0000FFF;
defparam prom_inst_12.INIT_RAM_06 = 256'hFFF0000FFC0007FFFFF00007FC0000000000001FF00007FFFFF0000FF80007FF;
defparam prom_inst_12.INIT_RAM_07 = 256'hFFF0000FFE0000000000001FF80007FFFFF0001FF80007FFFFE0000FFC0003FF;
defparam prom_inst_12.INIT_RAM_08 = 256'h0000003FF80003FFFFE0003FFC0003FFFFE0000FFC0003FFFFF0001FFE0003FF;
defparam prom_inst_12.INIT_RAM_09 = 256'hFFE0003FFE0003FFFFC0001FFE0001FFFFE0001FFE0001FFFFE0001FFE000000;
defparam prom_inst_12.INIT_RAM_0A = 256'hFFC0003FFF0000FFFFC0003FFF0001FFFFC0001FFF0000000000003FFC0003FF;
defparam prom_inst_12.INIT_RAM_0B = 256'hFFC0007FFF0000FFFFC0003FFF0000000000007FFE0001FFFFC0007FFE0001FF;
defparam prom_inst_12.INIT_RAM_0C = 256'hFF80003FFF800000000000FFFE0001FFFF80007FFF0001FFFF80003FFF0000FF;
defparam prom_inst_12.INIT_RAM_0D = 256'h000000FFFF0000FFFF8000FFFF0000FFFF00007FFF80007FFF80007FFF8000FF;
defparam prom_inst_12.INIT_RAM_0E = 256'hFF0001FFFF80007FFF0000FFFF80007FFF8000FFFFC0007FFF80007FFFC00000;
defparam prom_inst_12.INIT_RAM_0F = 256'hFE0000FFFFC0003FFF0000FFFFC0003FFF0000FFFFC00000000001FFFF00007F;
defparam prom_inst_12.INIT_RAM_10 = 256'hFE0001FFFFE0001FFE0000FFFFE00000000001FFFF80007FFF0001FFFF80007F;
defparam prom_inst_12.INIT_RAM_11 = 256'hFE0001FFFFE00000000003FFFFC0003FFE0003FFFFC0003FFE0001FFFFE0001F;
defparam prom_inst_12.INIT_RAM_12 = 256'h000007FFFFC0003FFC0003FFFFE0003FFC0001FFFFE0001FFE0003FFFFE0001F;
defparam prom_inst_12.INIT_RAM_13 = 256'hFC0007FFFFF0001FF80003FFFFF0000FFC0003FFFFF0000FFC0001FFFFF00000;
defparam prom_inst_12.INIT_RAM_14 = 256'hF80007FFFFF0000FFC0007FFFFF8000FFC0003FFFFF80000000007FFFFE0001F;
defparam prom_inst_12.INIT_RAM_15 = 256'hF8000FFFFFF80007F80007FFFFF8000000000FFFFFE0000FF8000FFFFFF0000F;
defparam prom_inst_12.INIT_RAM_16 = 256'hF00007FFFFFC000000000FFFFFF0000FF0000FFFFFF8000FF00007FFFFF80007;
defparam prom_inst_12.INIT_RAM_17 = 256'h00001FFFFFF80007F0001FFFFFF80007F0000FFFFFFC0003F0000FFFFFFC0003;
defparam prom_inst_12.INIT_RAM_18 = 256'hE0001FFFFFFC0007E0000FFFFFFC0003F0001FFFFFFC0003F0000FFFFFFC0000;
defparam prom_inst_12.INIT_RAM_19 = 256'hC0001FFFFFFE0001E0001FFFFFFE0001E0000FFFFFFE000000003FFFFFF80007;
defparam prom_inst_12.INIT_RAM_1A = 256'hE0003FFFFFFF0001E0001FFFFFFF000000003FFFFFFC0003E0003FFFFFFE0003;
defparam prom_inst_12.INIT_RAM_1B = 256'hC0003FFFFFFF000000007FFFFFFC0001C0007FFFFFFE0001C0003FFFFFFE0001;
defparam prom_inst_12.INIT_RAM_1C = 256'h0000FFFFFFFE000180007FFFFFFF000180003FFFFFFF0000C0007FFFFFFF0000;
defparam prom_inst_12.INIT_RAM_1D = 256'h8000FFFFFFFF000080007FFFFFFF800000007FFFFFFF800000003FFFFFFF8000;
defparam prom_inst_12.INIT_RAM_1E = 256'h00007FFFFFFF80000000FFFFFFFF800000007FFFFFFF80000000FFFFFFFF0000;
defparam prom_inst_12.INIT_RAM_1F = 256'h0000FFFFFFFFC00000007FFFFFFFC0000001FFFFFFFF00000000FFFFFFFF8000;
defparam prom_inst_12.INIT_RAM_20 = 256'h0000FFFFFFFFE0000001FFFFFFFF80000001FFFFFFFFC0000000FFFFFFFFC000;
defparam prom_inst_12.INIT_RAM_21 = 256'h0003FFFFFFFF80000003FFFFFFFFC0000001FFFFFFFFE0000001FFFFFFFFE000;
defparam prom_inst_12.INIT_RAM_22 = 256'h0003FFFFFFFFE0000001FFFFFFFFE0000003FFFFFFFFE0000001FFFFFFFFE000;
defparam prom_inst_12.INIT_RAM_23 = 256'h0003FFFFFFFFF0000003FFFFFFFFF0000001FFFFFFFFF0000007FFFFFFFFC000;
defparam prom_inst_12.INIT_RAM_24 = 256'h0007FFFFFFFFF0000003FFFFFFFFF0000007FFFFFFFFE0000007FFFFFFFFE000;
defparam prom_inst_12.INIT_RAM_25 = 256'h0003FFFFFFFFF800000FFFFFFFFFE0000007FFFFFFFFF0000007FFFFFFFFF000;
defparam prom_inst_12.INIT_RAM_26 = 256'h000FFFFFFFFFF000000FFFFFFFFFF8000007FFFFFFFFF8000007FFFFFFFFF800;
defparam prom_inst_12.INIT_RAM_27 = 256'h001FFFFFFFFFF800000FFFFFFFFFFC00000FFFFFFFFFFC000007FFFFFFFFFC00;
defparam prom_inst_12.INIT_RAM_28 = 256'h000FFFFFFFFFFC00001FFFFFFFFFFC00000FFFFFFFFFFC00001FFFFFFFFFF000;
defparam prom_inst_12.INIT_RAM_29 = 256'h001FFFFFFFFFFE00000FFFFFFFFFFC00003FFFFFFFFFF800001FFFFFFFFFFC00;
defparam prom_inst_12.INIT_RAM_2A = 256'h001FFFFFFFFFFC00003FFFFFFFFFFC00003FFFFFFFFFFC00001FFFFFFFFFFE00;
defparam prom_inst_12.INIT_RAM_2B = 256'h003FFFFFFFFFFC00003FFFFFFFFFFE00003FFFFFFFFFFE00003FFFFFFFFFFE00;
defparam prom_inst_12.INIT_RAM_2C = 256'h007FFFFFFFFFFE00003FFFFFFFFFFF00003FFFFFFFFFFF00001FFFFFFFFFF800;
defparam prom_inst_12.INIT_RAM_2D = 256'h007FFFFFFFFFFF00007FFFFFFFFFFF00003FFFFFFFFFF800003FFFFFFFFFFE00;
defparam prom_inst_12.INIT_RAM_2E = 256'h007FFFFFFFFFFF80003FFFFFFFFFF000001FFFFFFFFFFE00007FFFFFFFFFFF00;
defparam prom_inst_12.INIT_RAM_2F = 256'h007FFFFFFFFFF000000FFFFFFFFFFF0000FFFFFFFFFFFF80007FFFFFFFFFFF80;
defparam prom_inst_12.INIT_RAM_30 = 256'h000FFFFFFFFFFF80007FFFFFFFFFFF0000FFFFFFFFFFFFC0007FFFFFFFFFFF80;
defparam prom_inst_12.INIT_RAM_31 = 256'h007FFFFFFFFFFE0001FFFFFFFFFFFFC0003FFFFFFFFFFF0000FFFFFFFFFFE000;
defparam prom_inst_12.INIT_RAM_32 = 256'h01FFFFFFFFFFFFE0003FFFFFFFFFFE0000FFFFFFFFFFC0000007FFFFFFFFFF80;
defparam prom_inst_12.INIT_RAM_33 = 256'h001FFFFFFFFFFE0001FFFFFFFFFFC0000007FFFFFFFFFFC0003FFFFFFFFFFE00;
defparam prom_inst_12.INIT_RAM_34 = 256'h01FFFFFFFFFF80000003FFFFFFFFFFC0003FFFFFFFFFFC0003FFFFFFFFFFFFE0;
defparam prom_inst_12.INIT_RAM_35 = 256'h0001FFFFFFFFFFE0001FFFFFFFFFFC0003FFFFFFFFFFFFF0001FFFFFFFFFFC00;
defparam prom_inst_12.INIT_RAM_36 = 256'h000FFFFFFFFFF80007FFFFFFFFFFFFF8000FFFFFFFFFFC0003FFFFFFFFFF8000;
defparam prom_inst_12.INIT_RAM_37 = 256'h0FFFFFFFFFFFFFF80007FFFFFFFFF80007FFFFFFFFFF00000001FFFFFFFFFFF0;
defparam prom_inst_12.INIT_RAM_38 = 256'h0007FFFFFFFFF00007FFFFFFFFFE00000000FFFFFFFFFFF0000FFFFFFFFFF000;
defparam prom_inst_12.INIT_RAM_39 = 256'h0FFFFFFFFFFE00000000FFFFFFFFFFF80007FFFFFFFFF0000FFFFFFFFFFFFFFC;
defparam prom_inst_12.INIT_RAM_3A = 256'h00007FFFFFFFFFF80007FFFFFFFFE0001FFFFFFFFFFFFFFC0003FFFFFFFFF000;
defparam prom_inst_12.INIT_RAM_3B = 256'h0003FFFFFFFFE0001FFFFFFFFFFFFFFE0003FFFFFFFFE0000FFFFFFFFFFC0000;
defparam prom_inst_12.INIT_RAM_3C = 256'h3FFFFFFFFFFFFFFF0001FFFFFFFFE0001FFFFFFFFFFC000000003FFFFFFFFFFC;
defparam prom_inst_12.INIT_RAM_3D = 256'h0000FFFFFFFFC0003FFFFFFFFFF8000000003FFFFFFFFFFE0001FFFFFFFFC000;
defparam prom_inst_12.INIT_RAM_3E = 256'h3FFFFFFFFFF8000000001FFFFFFFFFFE0001FFFFFFFF80007FFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_3F = 256'h00001FFFFFFFFFFF0000FFFFFFFF80007FFFFFFFFFFFFFFF8000FFFFFFFF8000;

pROM prom_inst_13 (
    .DO({prom_inst_13_dout_w[30:0],prom_inst_13_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_11),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_13.READ_MODE = 1'b0;
defparam prom_inst_13.BIT_WIDTH = 1;
defparam prom_inst_13.RESET_MODE = "SYNC";
defparam prom_inst_13.INIT_RAM_00 = 256'h0000FFFFFFFF0000FFFFFFFFFFFFFFFF80007FFFFFFF80007FFFFFFFFFF00000;
defparam prom_inst_13.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFC0007FFFFFFF00007FFFFFFFFFE0000000000FFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_02 = 256'hE0003FFFFFFF0000FFFFFFFFFFE00000000007FFFFFFFFFF80007FFFFFFF0000;
defparam prom_inst_13.INIT_RAM_03 = 256'hFFFFFFFFFFC00000000007FFFFFFFFFFC0003FFFFFFE0001FFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_04 = 256'h000003FFFFFFFFFFC0003FFFFFFC0003FFFFFFFFFFFFFFFFE0001FFFFFFE0001;
defparam prom_inst_13.INIT_RAM_05 = 256'hE0001FFFFFFC0003FFFFFFFFFFFFFFFFF0001FFFFFFC0001FFFFFFFFFFC00000;
defparam prom_inst_13.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFF0000FFFFFFC0003FFFFFFFFFF800000000003FFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_07 = 256'hF8000FFFFFF80003FFFFFFFFFF000000000001FFFFFFFFFFE0001FFFFFF80007;
defparam prom_inst_13.INIT_RAM_08 = 256'hFFFFFFFFFF000000000000FFFFFFFFFFF0000FFFFFF80007FFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_09 = 256'h000000FFFFFFFFFFF00007FFFFF0000FFFFFFFFFFFFFFFFFFC0007FFFFF80007;
defparam prom_inst_13.INIT_RAM_0A = 256'hF80007FFFFE0001FFFFFFFFFFFFFFFFFFC0003FFFFF0000FFFFFFFFFFE000000;
defparam prom_inst_13.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFE0003FFFFE0000FFFFFFFFFFE0000000000007FFFFFFFFF;
defparam prom_inst_13.INIT_RAM_0C = 256'hFE0001FFFFE0001FFFFFFFFFFC0000000000007FFFFFFFFFFC0003FFFFE0001F;
defparam prom_inst_13.INIT_RAM_0D = 256'hFFFFFFFFF80000000000003FFFFFFFFFFC0003FFFFC0003FFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_0E = 256'h0000001FFFFFFFFFFE0001FFFF80003FFFFFFFFFFFFFFFFFFF0000FFFFC0001F;
defparam prom_inst_13.INIT_RAM_0F = 256'hFF0000FFFF80007FFFFFFFFFFFFFFFFFFF8000FFFFC0003FFFFFFFFFF8000000;
defparam prom_inst_13.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFFF80007FFF80003FFFFFFFFFF00000000000001FFFFFFFFF;
defparam prom_inst_13.INIT_RAM_11 = 256'hFFC0007FFF80007FFFFFFFFFF00000000000000FFFFFFFFFFF0000FFFF00007F;
defparam prom_inst_13.INIT_RAM_12 = 256'hFFFFFFFFE00000000000000FFFFFFFFFFF80007FFF0000FFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_13 = 256'h00000007FFFFFFFFFF80007FFE0001FFFFFFFFFFFFFFFFFFFFC0003FFF0000FF;
defparam prom_inst_13.INIT_RAM_14 = 256'hFFC0003FFE0001FFFFFFFFFFFFFFFFFFFFE0001FFE0001FFFFFFFFFFE0000000;
defparam prom_inst_13.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFE0001FFE0001FFFFFFFFFFC000000000000003FFFFFFFF;
defparam prom_inst_13.INIT_RAM_16 = 256'hFFF0000FFC0003FFFFFFFFFF8000000000000003FFFFFFFFFFE0003FFC0003FF;
defparam prom_inst_13.INIT_RAM_17 = 256'hFFFFFFFF8000000000000001FFFFFFFFFFE0001FF80003FFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_18 = 256'h00000001FFFFFFFFFFF0000FF80007FFFFFFFFFFFFFFFFFFFFF8000FFC0003FF;
defparam prom_inst_13.INIT_RAM_19 = 256'hFFF0000FF0000FFFFFFFFFFF7FFFFFFFFFF80007F80007FFFFFFFFFF00000000;
defparam prom_inst_13.INIT_RAM_1A = 256'hFFFFFFFE3FFFFFFFFFFC0003F0000FFFFFFFFFFF0000000000000000FFFFFFFF;
defparam prom_inst_13.INIT_RAM_1B = 256'hFFFC0003F0000FFFFFFFFFFE00000000000000007FFFFFFFFFF80007F0000FFF;
defparam prom_inst_13.INIT_RAM_1C = 256'hFFFFFFFC00000000000000007FFFFFFFFFFC0007E0001FFFFFFFFFFE3FFFFFFF;
defparam prom_inst_13.INIT_RAM_1D = 256'h000000003FFFFFFFFFFC0003C0001FFFFFFFFFFC1FFFFFFFFFFE0001E0001FFF;
defparam prom_inst_13.INIT_RAM_1E = 256'hFFFE0001C0003FFFFFFFFFF80FFFFFFFFFFF0001E0001FFFFFFFFFFC00000000;
defparam prom_inst_13.INIT_RAM_1F = 256'hFFFFFFF80FFFFFFFFFFF0000C0003FFFFFFFFFF800000000000000003FFFFFFF;
defparam prom_inst_13.INIT_RAM_20 = 256'hFFFF800080007FFFFFFFFFF800000000000000001FFFFFFFFFFE000180007FFF;
defparam prom_inst_13.INIT_RAM_21 = 256'hFFFFFFF000000000000000000FFFFFFFFFFF000080007FFFFFFFFFF007FFFFFF;
defparam prom_inst_13.INIT_RAM_22 = 256'h000000000FFFFFFFFFFF80000000FFFFFFFFFFF007FFFFFFFFFF800000007FFF;
defparam prom_inst_13.INIT_RAM_23 = 256'hFFFF80000001FFFFFFFFFFE003FFFFFFFFFFC0000000FFFFFFFFFFE000000000;
defparam prom_inst_13.INIT_RAM_24 = 256'hFFFFFFC001FFFFFFFFFFE0000000FFFFFFFFFFE0000000000000000007FFFFFF;
defparam prom_inst_13.INIT_RAM_25 = 256'hFFFFE0000001FFFFFFFFFFC0000000000000000003FFFFFFFFFFC0000001FFFF;
defparam prom_inst_13.INIT_RAM_26 = 256'hFFFFFF80000000000000000003FFFFFFFFFFC0000003FFFFFFFFFFC001FFFFFF;
defparam prom_inst_13.INIT_RAM_27 = 256'h0000000001FFFFFFFFFFE0000003FFFFFFFFFF8000FFFFFFFFFFF0000003FFFF;
defparam prom_inst_13.INIT_RAM_28 = 256'hFFFFF0000007FFFFFFFFFF8000FFFFFFFFFFF0000003FFFFFFFFFF8000000000;
defparam prom_inst_13.INIT_RAM_29 = 256'hFFFFFF00007FFFFFFFFFF8000007FFFFFFFFFF00000000000000000001FFFFFF;
defparam prom_inst_13.INIT_RAM_2A = 256'hFFFFFC000007FFFFFFFFFF00000000000000000000FFFFFFFFFFF000000FFFFF;
defparam prom_inst_13.INIT_RAM_2B = 256'hFFFFFE000000000000000000007FFFFFFFFFF800000FFFFFFFFFFE00003FFFFF;
defparam prom_inst_13.INIT_RAM_2C = 256'h00000000007FFFFFFFFFF800001FFFFFFFFFFE00003FFFFFFFFFFE00000FFFFF;
defparam prom_inst_13.INIT_RAM_2D = 256'hFFFFFC00003FFFFFFFFFFC00001FFFFFFFFFFE00001FFFFFFFFFFC0000000000;
defparam prom_inst_13.INIT_RAM_2E = 256'hFFFFFC00001FFFFFFFFFFF00001FFFFFFFFFFC000000000000000000003FFFFF;
defparam prom_inst_13.INIT_RAM_2F = 256'hFFFFFF00003FFFFFFFFFF8000000000000000000003FFFFFFFFFFE00003FFFFF;
defparam prom_inst_13.INIT_RAM_30 = 256'hFFFFF8000000000000000000001FFFFFFFFFFE00007FFFFFFFFFF800000FFFFF;
defparam prom_inst_13.INIT_RAM_31 = 256'h00000000000FFFFFFFFFFF00007FFFFFFFFFF0000007FFFFFFFFFF80003FFFFF;
defparam prom_inst_13.INIT_RAM_32 = 256'hFFFFFF0000FFFFFFFFFFF0000007FFFFFFFFFFC0007FFFFFFFFFF00000000000;
defparam prom_inst_13.INIT_RAM_33 = 256'hFFFFE0000003FFFFFFFFFFC000FFFFFFFFFFE0000000000000000000000FFFFF;
defparam prom_inst_13.INIT_RAM_34 = 256'hFFFFFFE000FFFFFFFFFFE00000000000000000000007FFFFFFFFFF8001FFFFFF;
defparam prom_inst_13.INIT_RAM_35 = 256'hFFFFC00000000000000000000007FFFFFFFFFFC001FFFFFFFFFFE0000003FFFF;
defparam prom_inst_13.INIT_RAM_36 = 256'h000000000003FFFFFFFFFFC003FFFFFFFFFFC0000001FFFFFFFFFFE001FFFFFF;
defparam prom_inst_13.INIT_RAM_37 = 256'hFFFFFFE003FFFFFFFFFFC0000001FFFFFFFFFFF001FFFFFFFFFFC00000000000;
defparam prom_inst_13.INIT_RAM_38 = 256'hFFFF80000000FFFFFFFFFFF003FFFFFFFFFF800000000000000000000003FFFF;
defparam prom_inst_13.INIT_RAM_39 = 256'hFFFFFFF803FFFFFFFFFF800000000000000000000001FFFFFFFFFFE007FFFFFF;
defparam prom_inst_13.INIT_RAM_3A = 256'hFFFF000000000000000000000000FFFFFFFFFFF007FFFFFFFFFF000000007FFF;
defparam prom_inst_13.INIT_RAM_3B = 256'h000000000000FFFFFFFFFFF00FFFFFFFFFFF000000007FFFFFFFFFFC07FFFFFF;
defparam prom_inst_13.INIT_RAM_3C = 256'hFFFFFFF81FFFFFFFFFFE000000003FFFFFFFFFFC0FFFFFFFFFFE000000000000;
defparam prom_inst_13.INIT_RAM_3D = 256'hFFFE000000001FFFFFFFFFFE0FFFFFFFFFFE0000000000000000000000007FFF;
defparam prom_inst_13.INIT_RAM_3E = 256'hFFFFFFFE1FFFFFFFFFFC0000000000000000000000007FFFFFFFFFFC1FFFFFFF;
defparam prom_inst_13.INIT_RAM_3F = 256'hFFFC0000000000000000000000003FFFFFFFFFFC3FFFFFFFFFFC000000001FFF;

pROM prom_inst_14 (
    .DO({prom_inst_14_dout_w[30:0],prom_inst_14_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_13),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_14.READ_MODE = 1'b0;
defparam prom_inst_14.BIT_WIDTH = 1;
defparam prom_inst_14.RESET_MODE = "SYNC";
defparam prom_inst_14.INIT_RAM_00 = 256'h0000000000001FFFFFFFFFFE3FFFFFFFFFF8000000000FFFFFFFFFFF1FFFFFFF;
defparam prom_inst_14.INIT_RAM_01 = 256'hFFFFFFFE7FFFFFFFFFF8000000000FFFFFFFFFFFBFFFFFFFFFF8000000000000;
defparam prom_inst_14.INIT_RAM_02 = 256'hFFF00000000007FFFFFFFFFFFFFFFFFFFFF80000000000000000000000001FFF;
defparam prom_inst_14.INIT_RAM_03 = 256'hFFFFFFFFFFFFFFFFFFF00000000000000000000000000FFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_04 = 256'hFFE00000000000000000000000000FFFFFFFFFFFFFFFFFFFFFE00000000003FF;
defparam prom_inst_14.INIT_RAM_05 = 256'h00000000000007FFFFFFFFFFFFFFFFFFFFE00000000003FFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFFFFC00000000001FFFFFFFFFFFFFFFFFFFFE0000000000000;
defparam prom_inst_14.INIT_RAM_07 = 256'hFFC00000000001FFFFFFFFFFFFFFFFFFFFC000000000000000000000000003FF;
defparam prom_inst_14.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFC000000000000000000000000003FFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_09 = 256'hFF8000000000000000000000000001FFFFFFFFFFFFFFFFFFFF800000000000FF;
defparam prom_inst_14.INIT_RAM_0A = 256'h00000000000001FFFFFFFFFFFFFFFFFFFF0000000000007FFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFF0000000000007FFFFFFFFFFFFFFFFFFF00000000000000;
defparam prom_inst_14.INIT_RAM_0C = 256'hFE0000000000003FFFFFFFFFFFFFFFFFFF0000000000000000000000000000FF;
defparam prom_inst_14.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFE00000000000000000000000000007FFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_0E = 256'hFE00000000000000000000000000007FFFFFFFFFFFFFFFFFFE0000000000003F;
defparam prom_inst_14.INIT_RAM_0F = 256'h000000000000003FFFFFFFFFFFFFFFFFFC0000000000001FFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFFFF80000000000000FFFFFFFFFFFFFFFFFFC00000000000000;
defparam prom_inst_14.INIT_RAM_11 = 256'hF80000000000000FFFFFFFFFFFFFFFFFF800000000000000000000000000003F;
defparam prom_inst_14.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFFFF800000000000000000000000000001FFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_13 = 256'hF000000000000000000000000000000FFFFFFFFFFFFFFFFFF000000000000007;
defparam prom_inst_14.INIT_RAM_14 = 256'h000000000000000FFFFFFFFFFFFFFFFFF000000000000007FFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFE000000000000003FFFFFFFFFFFFFFFFF000000000000000;
defparam prom_inst_14.INIT_RAM_16 = 256'hC000000000000001FFFFFFFFFFFFFFFFE0000000000000000000000000000007;
defparam prom_inst_14.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFC0000000000000000000000000000007FFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_18 = 256'hC0000000000000000000000000000003FFFFFFFFFFFFFFFFC000000000000001;
defparam prom_inst_14.INIT_RAM_19 = 256'h0000000000000001FFFFFFFFFFFFFFFF8000000000000000FFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFF8000000000000000FFFFFFFFFFFFFFFF8000000000000000;
defparam prom_inst_14.INIT_RAM_1B = 256'h00000000000000007FFFFFFFFFFFFFFF80000000000000000000000000000001;
defparam prom_inst_14.INIT_RAM_1C = 256'h3FFFFFFFFFFFFFFF00000000000000000000000000000000FFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_1D = 256'h00000000000000000000000000000000FFFFFFFFFFFFFFFE0000000000000000;
defparam prom_inst_14.INIT_RAM_1E = 256'h00000000000000007FFFFFFFFFFFFFFE00000000000000003FFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_1F = 256'h3FFFFFFFFFFFFFFC00000000000000001FFFFFFFFFFFFFFE0000000000000000;
defparam prom_inst_14.INIT_RAM_20 = 256'h00000000000000001FFFFFFFFFFFFFFC00000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_21 = 256'h0FFFFFFFFFFFFFFC000000000000000000000000000000003FFFFFFFFFFFFFFC;
defparam prom_inst_14.INIT_RAM_22 = 256'h000000000000000000000000000000001FFFFFFFFFFFFFF80000000000000000;
defparam prom_inst_14.INIT_RAM_23 = 256'h00000000000000001FFFFFFFFFFFFFF0000000000000000007FFFFFFFFFFFFF8;
defparam prom_inst_14.INIT_RAM_24 = 256'h0FFFFFFFFFFFFFF0000000000000000007FFFFFFFFFFFFF80000000000000000;
defparam prom_inst_14.INIT_RAM_25 = 256'h000000000000000003FFFFFFFFFFFFF000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_26 = 256'h03FFFFFFFFFFFFE00000000000000000000000000000000007FFFFFFFFFFFFE0;
defparam prom_inst_14.INIT_RAM_27 = 256'h0000000000000000000000000000000007FFFFFFFFFFFFE00000000000000000;
defparam prom_inst_14.INIT_RAM_28 = 256'h000000000000000003FFFFFFFFFFFFC0000000000000000001FFFFFFFFFFFFE0;
defparam prom_inst_14.INIT_RAM_29 = 256'h03FFFFFFFFFFFF80000000000000000001FFFFFFFFFFFFC00000000000000000;
defparam prom_inst_14.INIT_RAM_2A = 256'h000000000000000000FFFFFFFFFFFFC000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_2B = 256'h007FFFFFFFFFFF800000000000000000000000000000000001FFFFFFFFFFFF80;
defparam prom_inst_14.INIT_RAM_2C = 256'h0000000000000000000000000000000000FFFFFFFFFFFF000000000000000000;
defparam prom_inst_14.INIT_RAM_2D = 256'h000000000000000000FFFFFFFFFFFF000000000000000000007FFFFFFFFFFF00;
defparam prom_inst_14.INIT_RAM_2E = 256'h007FFFFFFFFFFE000000000000000000003FFFFFFFFFFF000000000000000000;
defparam prom_inst_14.INIT_RAM_2F = 256'h0000000000000000003FFFFFFFFFFE0000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_30 = 256'h001FFFFFFFFFFC0000000000000000000000000000000000003FFFFFFFFFFC00;
defparam prom_inst_14.INIT_RAM_31 = 256'h00000000000000000000000000000000003FFFFFFFFFFC000000000000000000;
defparam prom_inst_14.INIT_RAM_32 = 256'h0000000000000000001FFFFFFFFFF8000000000000000000000FFFFFFFFFFC00;
defparam prom_inst_14.INIT_RAM_33 = 256'h001FFFFFFFFFF8000000000000000000000FFFFFFFFFF8000000000000000000;
defparam prom_inst_14.INIT_RAM_34 = 256'h00000000000000000007FFFFFFFFF80000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_35 = 256'h0007FFFFFFFFF00000000000000000000000000000000000000FFFFFFFFFF000;
defparam prom_inst_14.INIT_RAM_36 = 256'h000000000000000000000000000000000007FFFFFFFFE0000000000000000000;
defparam prom_inst_14.INIT_RAM_37 = 256'h00000000000000000007FFFFFFFFE00000000000000000000003FFFFFFFFE000;
defparam prom_inst_14.INIT_RAM_38 = 256'h0003FFFFFFFFC00000000000000000000001FFFFFFFFE0000000000000000000;
defparam prom_inst_14.INIT_RAM_39 = 256'h00000000000000000001FFFFFFFFC00000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_3A = 256'h0000FFFFFFFFC000000000000000000000000000000000000003FFFFFFFFC000;
defparam prom_inst_14.INIT_RAM_3B = 256'h000000000000000000000000000000000001FFFFFFFF80000000000000000000;
defparam prom_inst_14.INIT_RAM_3C = 256'h00000000000000000000FFFFFFFF000000000000000000000000FFFFFFFF8000;
defparam prom_inst_14.INIT_RAM_3D = 256'h0000FFFFFFFF0000000000000000000000007FFFFFFF80000000000000000000;
defparam prom_inst_14.INIT_RAM_3E = 256'h000000000000000000003FFFFFFF000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_3F = 256'h00003FFFFFFE00000000000000000000000000000000000000007FFFFFFE0000;

pROM prom_inst_15 (
    .DO({prom_inst_15_dout_w[30:0],prom_inst_15_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_15),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_15.READ_MODE = 1'b0;
defparam prom_inst_15.BIT_WIDTH = 1;
defparam prom_inst_15.RESET_MODE = "SYNC";
defparam prom_inst_15.INIT_RAM_00 = 256'h0000000000000000000000000000000000007FFFFFFE00000000000000000000;
defparam prom_inst_15.INIT_RAM_01 = 256'h000000000000000000003FFFFFFC0000000000000000000000001FFFFFFE0000;
defparam prom_inst_15.INIT_RAM_02 = 256'h00003FFFFFFC0000000000000000000000001FFFFFFC00000000000000000000;
defparam prom_inst_15.INIT_RAM_03 = 256'h000000000000000000000FFFFFFC000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_04 = 256'h000007FFFFF800000000000000000000000000000000000000001FFFFFF80000;
defparam prom_inst_15.INIT_RAM_05 = 256'h0000000000000000000000000000000000000FFFFFF000000000000000000000;
defparam prom_inst_15.INIT_RAM_06 = 256'h000000000000000000000FFFFFF000000000000000000000000007FFFFF80000;
defparam prom_inst_15.INIT_RAM_07 = 256'h000007FFFFE000000000000000000000000003FFFFF000000000000000000000;
defparam prom_inst_15.INIT_RAM_08 = 256'h0000000000000000000001FFFFE0000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_09 = 256'h000001FFFFE0000000000000000000000000000000000000000007FFFFC00000;
defparam prom_inst_15.INIT_RAM_0A = 256'h00000000000000000000000000000000000003FFFFC000000000000000000000;
defparam prom_inst_15.INIT_RAM_0B = 256'h0000000000000000000001FFFF8000000000000000000000000000FFFFC00000;
defparam prom_inst_15.INIT_RAM_0C = 256'h000001FFFF8000000000000000000000000000FFFFC000000000000000000000;
defparam prom_inst_15.INIT_RAM_0D = 256'h00000000000000000000007FFF80000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_0E = 256'h0000003FFF00000000000000000000000000000000000000000000FFFF000000;
defparam prom_inst_15.INIT_RAM_0F = 256'h00000000000000000000000000000000000000FFFE0000000000000000000000;
defparam prom_inst_15.INIT_RAM_10 = 256'h00000000000000000000007FFE00000000000000000000000000003FFF000000;
defparam prom_inst_15.INIT_RAM_11 = 256'h0000003FFC00000000000000000000000000001FFE0000000000000000000000;
defparam prom_inst_15.INIT_RAM_12 = 256'h00000000000000000000001FFE00000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_13 = 256'h0000000FFC000000000000000000000000000000000000000000003FFC000000;
defparam prom_inst_15.INIT_RAM_14 = 256'h000000000000000000000000000000000000001FF80000000000000000000000;
defparam prom_inst_15.INIT_RAM_15 = 256'h00000000000000000000001FF0000000000000000000000000000007F8000000;
defparam prom_inst_15.INIT_RAM_16 = 256'h0000000FF0000000000000000000000000000007F80000000000000000000000;
defparam prom_inst_15.INIT_RAM_17 = 256'h000000000000000000000003F000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_18 = 256'h00000003F00000000000000000000000000000000000000000000007E0000000;
defparam prom_inst_15.INIT_RAM_19 = 256'h0000000000000000000000000000000000000007E00000000000000000000000;
defparam prom_inst_15.INIT_RAM_1A = 256'h000000000000000000000003C0000000000000000000000000000001E0000000;
defparam prom_inst_15.INIT_RAM_1B = 256'h0000000380000000000000000000000000000000C00000000000000000000000;
defparam prom_inst_15.INIT_RAM_1C = 256'h000000000000000000000000C000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000180000000;
defparam prom_inst_15.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_16 (
    .DO({prom_inst_16_dout_w[30:0],prom_inst_16_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_17),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_16.READ_MODE = 1'b0;
defparam prom_inst_16.BIT_WIDTH = 1;
defparam prom_inst_16.RESET_MODE = "SYNC";
defparam prom_inst_16.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_16.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_17 (
    .DO({prom_inst_17_dout_w[30:0],prom_inst_17_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_17),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_17.READ_MODE = 1'b0;
defparam prom_inst_17.BIT_WIDTH = 1;
defparam prom_inst_17.RESET_MODE = "SYNC";
defparam prom_inst_17.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_17.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_18 (
    .DO({prom_inst_18_dout_w[29:0],prom_inst_18_dout[1:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_19),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_18.READ_MODE = 1'b0;
defparam prom_inst_18.BIT_WIDTH = 2;
defparam prom_inst_18.RESET_MODE = "SYNC";
defparam prom_inst_18.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_18.INIT_RAM_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[17]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(ad[16]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(ad[15]),
  .CLK(clk),
  .CE(ce)
);
DFFE dff_inst_3 (
  .Q(dff_q_3),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce)
);
MUX2 mux_inst_10 (
  .O(mux_o_10),
  .I0(prom_inst_0_dout[0]),
  .I1(prom_inst_1_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_11 (
  .O(mux_o_11),
  .I0(prom_inst_2_dout[0]),
  .I1(prom_inst_3_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_12 (
  .O(mux_o_12),
  .I0(prom_inst_4_dout[0]),
  .I1(prom_inst_5_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_13 (
  .O(mux_o_13),
  .I0(prom_inst_6_dout[0]),
  .I1(prom_inst_7_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_14 (
  .O(mux_o_14),
  .I0(prom_inst_16_dout[0]),
  .I1(prom_inst_18_dout[0]),
  .S0(dff_q_3)
);
MUX2 mux_inst_15 (
  .O(mux_o_15),
  .I0(mux_o_10),
  .I1(mux_o_11),
  .S0(dff_q_2)
);
MUX2 mux_inst_16 (
  .O(mux_o_16),
  .I0(mux_o_12),
  .I1(mux_o_13),
  .S0(dff_q_2)
);
MUX2 mux_inst_18 (
  .O(mux_o_18),
  .I0(mux_o_15),
  .I1(mux_o_16),
  .S0(dff_q_1)
);
MUX2 mux_inst_20 (
  .O(dout[0]),
  .I0(mux_o_18),
  .I1(mux_o_14),
  .S0(dff_q_0)
);
MUX2 mux_inst_31 (
  .O(mux_o_31),
  .I0(prom_inst_8_dout[1]),
  .I1(prom_inst_9_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_32 (
  .O(mux_o_32),
  .I0(prom_inst_10_dout[1]),
  .I1(prom_inst_11_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_33 (
  .O(mux_o_33),
  .I0(prom_inst_12_dout[1]),
  .I1(prom_inst_13_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_34 (
  .O(mux_o_34),
  .I0(prom_inst_14_dout[1]),
  .I1(prom_inst_15_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_35 (
  .O(mux_o_35),
  .I0(prom_inst_17_dout[1]),
  .I1(prom_inst_18_dout[1]),
  .S0(dff_q_3)
);
MUX2 mux_inst_36 (
  .O(mux_o_36),
  .I0(mux_o_31),
  .I1(mux_o_32),
  .S0(dff_q_2)
);
MUX2 mux_inst_37 (
  .O(mux_o_37),
  .I0(mux_o_33),
  .I1(mux_o_34),
  .S0(dff_q_2)
);
MUX2 mux_inst_39 (
  .O(mux_o_39),
  .I0(mux_o_36),
  .I1(mux_o_37),
  .S0(dff_q_1)
);
MUX2 mux_inst_41 (
  .O(dout[1]),
  .I0(mux_o_39),
  .I1(mux_o_35),
  .S0(dff_q_0)
);
endmodule //Gowin_pROM
